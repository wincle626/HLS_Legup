// legup_system.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module legup_system (
		input  wire        clk_clk,                      //                    clk.clk
		input  wire [2:0]  leap_debug_port_select,       //        leap_debug_port.select
		output wire [17:0] leap_debug_port_lights,       //                       .lights
		output wire        leap_profiling_signals_start, // leap_profiling_signals.start
		output wire        leap_profiling_signals_end,   //                       .end
		input  wire        reset_reset_n,                //                  reset.reset_n
		output wire [12:0] sdram_wire_addr,              //             sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                //                       .ba
		output wire        sdram_wire_cas_n,             //                       .cas_n
		output wire        sdram_wire_cke,               //                       .cke
		output wire        sdram_wire_cs_n,              //                       .cs_n
		inout  wire [15:0] sdram_wire_dq,                //                       .dq
		output wire [1:0]  sdram_wire_dqm,               //                       .dqm
		output wire        sdram_wire_ras_n,             //                       .ras_n
		output wire        sdram_wire_we_n               //                       .we_n
	);

	wire  [31:0] tiger_mips_instruction_master_readdata;                    // Leap_Profiler:avs_from_cpu_readdata -> Tiger_MIPS:avm_instrMaster_readdata
	wire         tiger_mips_instruction_master_waitrequest;                 // Leap_Profiler:avs_from_cpu_waitrequest -> Tiger_MIPS:avm_instrMaster_waitrequest
	wire  [31:0] tiger_mips_instruction_master_address;                     // Tiger_MIPS:avm_instrMaster_address -> Leap_Profiler:avs_from_cpu_address
	wire         tiger_mips_instruction_master_read;                        // Tiger_MIPS:avm_instrMaster_read -> Leap_Profiler:avs_from_cpu_read
	wire   [3:0] tiger_mips_instruction_master_byteenable;                  // Tiger_MIPS:avm_instrMaster_byteenable -> Leap_Profiler:avs_from_cpu_byteenable
	wire         tiger_mips_instruction_master_readdatavalid;               // Leap_Profiler:avs_from_cpu_readdatavalid -> Tiger_MIPS:avm_instrMaster_readdatavalid
	wire         tiger_mips_instruction_master_write;                       // Tiger_MIPS:avm_instrMaster_write -> Leap_Profiler:avs_from_cpu_write
	wire  [31:0] tiger_mips_instruction_master_writedata;                   // Tiger_MIPS:avm_instrMaster_writedata -> Leap_Profiler:avs_from_cpu_writedata
	wire  [31:0] leap_sim_control_bridge_master_readdata;                   // mm_interconnect_0:Leap_Sim_Control_bridge_master_readdata -> Leap_Sim_Control:avm_bridge_master_readdata
	wire         leap_sim_control_bridge_master_waitrequest;                // mm_interconnect_0:Leap_Sim_Control_bridge_master_waitrequest -> Leap_Sim_Control:avm_bridge_master_waitrequest
	wire  [31:0] leap_sim_control_bridge_master_address;                    // Leap_Sim_Control:avm_bridge_master_address -> mm_interconnect_0:Leap_Sim_Control_bridge_master_address
	wire   [3:0] leap_sim_control_bridge_master_byteenable;                 // Leap_Sim_Control:avm_bridge_master_byteenable -> mm_interconnect_0:Leap_Sim_Control_bridge_master_byteenable
	wire         leap_sim_control_bridge_master_read;                       // Leap_Sim_Control:avm_bridge_master_read -> mm_interconnect_0:Leap_Sim_Control_bridge_master_read
	wire         leap_sim_control_bridge_master_write;                      // Leap_Sim_Control:avm_bridge_master_write -> mm_interconnect_0:Leap_Sim_Control_bridge_master_write
	wire  [31:0] leap_sim_control_bridge_master_writedata;                  // Leap_Sim_Control:avm_bridge_master_writedata -> mm_interconnect_0:Leap_Sim_Control_bridge_master_writedata
	wire  [31:0] mm_interconnect_0_leap_profiler_leapslave_readdata;        // Leap_Profiler:avs_leapSlave_readdata -> mm_interconnect_0:Leap_Profiler_leapslave_readdata
	wire  [29:0] mm_interconnect_0_leap_profiler_leapslave_address;         // mm_interconnect_0:Leap_Profiler_leapslave_address -> Leap_Profiler:avs_leapSlave_address
	wire         mm_interconnect_0_leap_profiler_leapslave_read;            // mm_interconnect_0:Leap_Profiler_leapslave_read -> Leap_Profiler:avs_leapSlave_read
	wire         mm_interconnect_0_leap_profiler_leapslave_write;           // mm_interconnect_0:Leap_Profiler_leapslave_write -> Leap_Profiler:avs_leapSlave_write
	wire  [31:0] mm_interconnect_0_leap_profiler_leapslave_writedata;       // mm_interconnect_0:Leap_Profiler_leapslave_writedata -> Leap_Profiler:avs_leapSlave_writedata
	wire  [31:0] dcache_cache_master_readdata;                              // mm_interconnect_1:DCache_cache_master_readdata -> DCache:avm_cache_readdata
	wire         dcache_cache_master_waitrequest;                           // mm_interconnect_1:DCache_cache_master_waitrequest -> DCache:avm_cache_waitrequest
	wire  [31:0] dcache_cache_master_address;                               // DCache:avm_cache_address -> mm_interconnect_1:DCache_cache_master_address
	wire   [3:0] dcache_cache_master_byteenable;                            // DCache:avm_cache_byteenable -> mm_interconnect_1:DCache_cache_master_byteenable
	wire         dcache_cache_master_read;                                  // DCache:avm_cache_read -> mm_interconnect_1:DCache_cache_master_read
	wire         dcache_cache_master_readdatavalid;                         // mm_interconnect_1:DCache_cache_master_readdatavalid -> DCache:avm_cache_readdatavalid
	wire         dcache_cache_master_write;                                 // DCache:avm_cache_write -> mm_interconnect_1:DCache_cache_master_write
	wire  [31:0] dcache_cache_master_writedata;                             // DCache:avm_cache_writedata -> mm_interconnect_1:DCache_cache_master_writedata
	wire   [2:0] dcache_cache_master_burstcount;                            // DCache:avm_cache_burstcount -> mm_interconnect_1:DCache_cache_master_burstcount
	wire         tiger_icache_icache_master_beginbursttransfer;             // Tiger_ICache:avm_icache_master_beginbursttransfer -> mm_interconnect_1:Tiger_ICache_icache_master_beginbursttransfer
	wire  [31:0] tiger_icache_icache_master_readdata;                       // mm_interconnect_1:Tiger_ICache_icache_master_readdata -> Tiger_ICache:avm_icache_master_readdata
	wire         tiger_icache_icache_master_waitrequest;                    // mm_interconnect_1:Tiger_ICache_icache_master_waitrequest -> Tiger_ICache:avm_icache_master_waitrequest
	wire  [31:0] tiger_icache_icache_master_address;                        // Tiger_ICache:avm_icache_master_address -> mm_interconnect_1:Tiger_ICache_icache_master_address
	wire         tiger_icache_icache_master_read;                           // Tiger_ICache:avm_icache_master_read -> mm_interconnect_1:Tiger_ICache_icache_master_read
	wire         tiger_icache_icache_master_readdatavalid;                  // mm_interconnect_1:Tiger_ICache_icache_master_readdatavalid -> Tiger_ICache:avm_icache_master_readdatavalid
	wire   [5:0] tiger_icache_icache_master_burstcount;                     // Tiger_ICache:avm_icache_master_burstcount -> mm_interconnect_1:Tiger_ICache_icache_master_burstcount
	wire  [31:0] jtag_to_fpga_bridge_master_readdata;                       // mm_interconnect_1:JTAG_to_FPGA_Bridge_master_readdata -> JTAG_to_FPGA_Bridge:master_readdata
	wire         jtag_to_fpga_bridge_master_waitrequest;                    // mm_interconnect_1:JTAG_to_FPGA_Bridge_master_waitrequest -> JTAG_to_FPGA_Bridge:master_waitrequest
	wire  [31:0] jtag_to_fpga_bridge_master_address;                        // JTAG_to_FPGA_Bridge:master_address -> mm_interconnect_1:JTAG_to_FPGA_Bridge_master_address
	wire         jtag_to_fpga_bridge_master_read;                           // JTAG_to_FPGA_Bridge:master_read -> mm_interconnect_1:JTAG_to_FPGA_Bridge_master_read
	wire   [3:0] jtag_to_fpga_bridge_master_byteenable;                     // JTAG_to_FPGA_Bridge:master_byteenable -> mm_interconnect_1:JTAG_to_FPGA_Bridge_master_byteenable
	wire         jtag_to_fpga_bridge_master_readdatavalid;                  // mm_interconnect_1:JTAG_to_FPGA_Bridge_master_readdatavalid -> JTAG_to_FPGA_Bridge:master_readdatavalid
	wire         jtag_to_fpga_bridge_master_write;                          // JTAG_to_FPGA_Bridge:master_write -> mm_interconnect_1:JTAG_to_FPGA_Bridge_master_write
	wire  [31:0] jtag_to_fpga_bridge_master_writedata;                      // JTAG_to_FPGA_Bridge:master_writedata -> mm_interconnect_1:JTAG_to_FPGA_Bridge_master_writedata
	wire  [31:0] tiger_mips_data_master_readdata;                           // mm_interconnect_1:Tiger_MIPS_data_master_readdata -> Tiger_MIPS:avm_dataMaster_readdata
	wire         tiger_mips_data_master_waitrequest;                        // mm_interconnect_1:Tiger_MIPS_data_master_waitrequest -> Tiger_MIPS:avm_dataMaster_waitrequest
	wire  [31:0] tiger_mips_data_master_address;                            // Tiger_MIPS:avm_dataMaster_address -> mm_interconnect_1:Tiger_MIPS_data_master_address
	wire         tiger_mips_data_master_read;                               // Tiger_MIPS:avm_dataMaster_read -> mm_interconnect_1:Tiger_MIPS_data_master_read
	wire   [3:0] tiger_mips_data_master_byteenable;                         // Tiger_MIPS:avm_dataMaster_byteenable -> mm_interconnect_1:Tiger_MIPS_data_master_byteenable
	wire         tiger_mips_data_master_readdatavalid;                      // mm_interconnect_1:Tiger_MIPS_data_master_readdatavalid -> Tiger_MIPS:avm_dataMaster_readdatavalid
	wire         tiger_mips_data_master_write;                              // Tiger_MIPS:avm_dataMaster_write -> mm_interconnect_1:Tiger_MIPS_data_master_write
	wire  [31:0] tiger_mips_data_master_writedata;                          // Tiger_MIPS:avm_dataMaster_writedata -> mm_interconnect_1:Tiger_MIPS_data_master_writedata
	wire         mm_interconnect_1_sdram_s1_chipselect;                     // mm_interconnect_1:SDRAM_s1_chipselect -> SDRAM:az_cs
	wire  [15:0] mm_interconnect_1_sdram_s1_readdata;                       // SDRAM:za_data -> mm_interconnect_1:SDRAM_s1_readdata
	wire         mm_interconnect_1_sdram_s1_waitrequest;                    // SDRAM:za_waitrequest -> mm_interconnect_1:SDRAM_s1_waitrequest
	wire  [24:0] mm_interconnect_1_sdram_s1_address;                        // mm_interconnect_1:SDRAM_s1_address -> SDRAM:az_addr
	wire         mm_interconnect_1_sdram_s1_read;                           // mm_interconnect_1:SDRAM_s1_read -> SDRAM:az_rd_n
	wire   [1:0] mm_interconnect_1_sdram_s1_byteenable;                     // mm_interconnect_1:SDRAM_s1_byteenable -> SDRAM:az_be_n
	wire         mm_interconnect_1_sdram_s1_readdatavalid;                  // SDRAM:za_valid -> mm_interconnect_1:SDRAM_s1_readdatavalid
	wire         mm_interconnect_1_sdram_s1_write;                          // mm_interconnect_1:SDRAM_s1_write -> SDRAM:az_wr_n
	wire  [15:0] mm_interconnect_1_sdram_s1_writedata;                      // mm_interconnect_1:SDRAM_s1_writedata -> SDRAM:az_data
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_1:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;    // JTAG_UART:av_readdata -> mm_interconnect_1:JTAG_UART_avalon_jtag_slave_readdata
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest; // JTAG_UART:av_waitrequest -> mm_interconnect_1:JTAG_UART_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_1:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_1:JTAG_UART_avalon_jtag_slave_read -> JTAG_UART:av_read_n
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_1:JTAG_UART_avalon_jtag_slave_write -> JTAG_UART:av_write_n
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_1:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	wire  [31:0] mm_interconnect_1_leap_sim_control_bridge_slave_readdata;  // Leap_Sim_Control:avs_bridge_slave_readdata -> mm_interconnect_1:Leap_Sim_Control_bridge_slave_readdata
	wire   [7:0] mm_interconnect_1_leap_sim_control_bridge_slave_address;   // mm_interconnect_1:Leap_Sim_Control_bridge_slave_address -> Leap_Sim_Control:avs_bridge_slave_address
	wire         mm_interconnect_1_leap_sim_control_bridge_slave_read;      // mm_interconnect_1:Leap_Sim_Control_bridge_slave_read -> Leap_Sim_Control:avs_bridge_slave_read
	wire         mm_interconnect_1_leap_sim_control_bridge_slave_write;     // mm_interconnect_1:Leap_Sim_Control_bridge_slave_write -> Leap_Sim_Control:avs_bridge_slave_write
	wire  [31:0] mm_interconnect_1_leap_sim_control_bridge_slave_writedata; // mm_interconnect_1:Leap_Sim_Control_bridge_slave_writedata -> Leap_Sim_Control:avs_bridge_slave_writedata
	wire  [31:0] mm_interconnect_1_dcache_cache_slave_readdata;             // DCache:avs_cache_readdata -> mm_interconnect_1:DCache_cache_slave_readdata
	wire         mm_interconnect_1_dcache_cache_slave_waitrequest;          // DCache:avs_cache_waitrequest -> mm_interconnect_1:DCache_cache_slave_waitrequest
	wire  [30:0] mm_interconnect_1_dcache_cache_slave_address;              // mm_interconnect_1:DCache_cache_slave_address -> DCache:avs_cache_address
	wire         mm_interconnect_1_dcache_cache_slave_read;                 // mm_interconnect_1:DCache_cache_slave_read -> DCache:avs_cache_read
	wire   [3:0] mm_interconnect_1_dcache_cache_slave_byteenable;           // mm_interconnect_1:DCache_cache_slave_byteenable -> DCache:avs_cache_byteenable
	wire         mm_interconnect_1_dcache_cache_slave_readdatavalid;        // DCache:avs_cache_readdatavalid -> mm_interconnect_1:DCache_cache_slave_readdatavalid
	wire         mm_interconnect_1_dcache_cache_slave_write;                // mm_interconnect_1:DCache_cache_slave_write -> DCache:avs_cache_write
	wire  [31:0] mm_interconnect_1_dcache_cache_slave_writedata;            // mm_interconnect_1:DCache_cache_slave_writedata -> DCache:avs_cache_writedata
	wire  [31:0] leap_profiler_to_memory_readdata;                          // mm_interconnect_3:Leap_Profiler_to_memory_readdata -> Leap_Profiler:avs_to_memory_readdata
	wire         leap_profiler_to_memory_waitrequest;                       // mm_interconnect_3:Leap_Profiler_to_memory_waitrequest -> Leap_Profiler:avs_to_memory_waitrequest
	wire  [31:0] leap_profiler_to_memory_address;                           // Leap_Profiler:avs_to_memory_address -> mm_interconnect_3:Leap_Profiler_to_memory_address
	wire         leap_profiler_to_memory_read;                              // Leap_Profiler:avs_to_memory_read -> mm_interconnect_3:Leap_Profiler_to_memory_read
	wire   [3:0] leap_profiler_to_memory_byteenable;                        // Leap_Profiler:avs_to_memory_byteenable -> mm_interconnect_3:Leap_Profiler_to_memory_byteenable
	wire         leap_profiler_to_memory_readdatavalid;                     // mm_interconnect_3:Leap_Profiler_to_memory_readdatavalid -> Leap_Profiler:avs_to_memory_readdatavalid
	wire         leap_profiler_to_memory_write;                             // Leap_Profiler:avs_to_memory_write -> mm_interconnect_3:Leap_Profiler_to_memory_write
	wire  [31:0] leap_profiler_to_memory_writedata;                         // Leap_Profiler:avs_to_memory_writedata -> mm_interconnect_3:Leap_Profiler_to_memory_writedata
	wire  [31:0] mm_interconnect_3_tiger_icache_icache_slave_readdata;      // Tiger_ICache:avs_icache_slave_readdata -> mm_interconnect_3:Tiger_ICache_icache_slave_readdata
	wire         mm_interconnect_3_tiger_icache_icache_slave_waitrequest;   // Tiger_ICache:avs_icache_slave_waitrequest -> mm_interconnect_3:Tiger_ICache_icache_slave_waitrequest
	wire  [29:0] mm_interconnect_3_tiger_icache_icache_slave_address;       // mm_interconnect_3:Tiger_ICache_icache_slave_address -> Tiger_ICache:avs_icache_slave_address
	wire         mm_interconnect_3_tiger_icache_icache_slave_read;          // mm_interconnect_3:Tiger_ICache_icache_slave_read -> Tiger_ICache:avs_icache_slave_read
	wire         mm_interconnect_3_tiger_icache_icache_slave_readdatavalid; // Tiger_ICache:avs_icache_slave_readdatavalid -> mm_interconnect_3:Tiger_ICache_icache_slave_readdatavalid
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [DCache:reset, JTAG_UART:rst_n, Leap_Profiler:reset, Leap_Sim_Control:reset, SDRAM:reset_n, Tiger_ICache:reset_n, mm_interconnect_0:Leap_Sim_Control_reset_reset_bridge_in_reset_reset, mm_interconnect_1:DCache_reset_reset_bridge_in_reset_reset, mm_interconnect_1:JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_3:Leap_Profiler_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [Tiger_MIPS:reset, mm_interconnect_1:Tiger_MIPS_reset_reset_bridge_in_reset_reset]
	wire         leap_profiler_leap_processor_reset_reset;                  // Leap_Profiler:tiger_soft_reset -> rst_controller_001:reset_in1

	legup_dm_wt_cache dcache (
		.reset                   (rst_controller_reset_out_reset),                     //        reset.reset
		.clk                     (clk_clk),                                            //          clk.clk
		.avs_cache_address       (mm_interconnect_1_dcache_cache_slave_address),       //  cache_slave.address
		.avs_cache_byteenable    (mm_interconnect_1_dcache_cache_slave_byteenable),    //             .byteenable
		.avs_cache_read          (mm_interconnect_1_dcache_cache_slave_read),          //             .read
		.avs_cache_write         (mm_interconnect_1_dcache_cache_slave_write),         //             .write
		.avs_cache_writedata     (mm_interconnect_1_dcache_cache_slave_writedata),     //             .writedata
		.avs_cache_readdata      (mm_interconnect_1_dcache_cache_slave_readdata),      //             .readdata
		.avs_cache_readdatavalid (mm_interconnect_1_dcache_cache_slave_readdatavalid), //             .readdatavalid
		.avs_cache_waitrequest   (mm_interconnect_1_dcache_cache_slave_waitrequest),   //             .waitrequest
		.avm_cache_readdata      (dcache_cache_master_readdata),                       // cache_master.readdata
		.avm_cache_readdatavalid (dcache_cache_master_readdatavalid),                  //             .readdatavalid
		.avm_cache_waitrequest   (dcache_cache_master_waitrequest),                    //             .waitrequest
		.avm_cache_address       (dcache_cache_master_address),                        //             .address
		.avm_cache_burstcount    (dcache_cache_master_burstcount),                     //             .burstcount
		.avm_cache_byteenable    (dcache_cache_master_byteenable),                     //             .byteenable
		.avm_cache_read          (dcache_cache_master_read),                           //             .read
		.avm_cache_write         (dcache_cache_master_write),                          //             .write
		.avm_cache_writedata     (dcache_cache_master_writedata)                       //             .writedata
	);

	legup_system_JTAG_UART jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         ()                                                           //               irq.irq
	);

	legup_system_JTAG_to_FPGA_Bridge #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) jtag_to_fpga_bridge (
		.clk_clk              (clk_clk),                                  //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                           //    clk_reset.reset
		.master_address       (jtag_to_fpga_bridge_master_address),       //       master.address
		.master_readdata      (jtag_to_fpga_bridge_master_readdata),      //             .readdata
		.master_read          (jtag_to_fpga_bridge_master_read),          //             .read
		.master_write         (jtag_to_fpga_bridge_master_write),         //             .write
		.master_writedata     (jtag_to_fpga_bridge_master_writedata),     //             .writedata
		.master_waitrequest   (jtag_to_fpga_bridge_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (jtag_to_fpga_bridge_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (jtag_to_fpga_bridge_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                          // master_reset.reset
	);

	LeapTop #(
		.STARTING_PC   (1073741856),
		.prof_param_N2 (8),
		.prof_param_S2 (5),
		.prof_param_CW (32)
	) leap_profiler (
		.clk                         (clk_clk),                                             //                clock.clk
		.reset                       (rst_controller_reset_out_reset),                      //                reset.reset
		.tiger_soft_reset            (leap_profiler_leap_processor_reset_reset),            // leap_processor_reset.reset
		.avs_from_cpu_address        (tiger_mips_instruction_master_address),               //             from_cpu.address
		.avs_from_cpu_read           (tiger_mips_instruction_master_read),                  //                     .read
		.avs_from_cpu_write          (tiger_mips_instruction_master_write),                 //                     .write
		.avs_from_cpu_writedata      (tiger_mips_instruction_master_writedata),             //                     .writedata
		.avs_from_cpu_byteenable     (tiger_mips_instruction_master_byteenable),            //                     .byteenable
		.avs_from_cpu_readdata       (tiger_mips_instruction_master_readdata),              //                     .readdata
		.avs_from_cpu_waitrequest    (tiger_mips_instruction_master_waitrequest),           //                     .waitrequest
		.avs_from_cpu_readdatavalid  (tiger_mips_instruction_master_readdatavalid),         //                     .readdatavalid
		.avs_to_memory_address       (leap_profiler_to_memory_address),                     //            to_memory.address
		.avs_to_memory_read          (leap_profiler_to_memory_read),                        //                     .read
		.avs_to_memory_write         (leap_profiler_to_memory_write),                       //                     .write
		.avs_to_memory_writedata     (leap_profiler_to_memory_writedata),                   //                     .writedata
		.avs_to_memory_byteenable    (leap_profiler_to_memory_byteenable),                  //                     .byteenable
		.avs_to_memory_readdata      (leap_profiler_to_memory_readdata),                    //                     .readdata
		.avs_to_memory_waitrequest   (leap_profiler_to_memory_waitrequest),                 //                     .waitrequest
		.avs_to_memory_readdatavalid (leap_profiler_to_memory_readdatavalid),               //                     .readdatavalid
		.avs_leapSlave_address       (mm_interconnect_0_leap_profiler_leapslave_address),   //            leapslave.address
		.avs_leapSlave_read          (mm_interconnect_0_leap_profiler_leapslave_read),      //                     .read
		.avs_leapSlave_write         (mm_interconnect_0_leap_profiler_leapslave_write),     //                     .write
		.avs_leapSlave_writedata     (mm_interconnect_0_leap_profiler_leapslave_writedata), //                     .writedata
		.avs_leapSlave_readdata      (mm_interconnect_0_leap_profiler_leapslave_readdata),  //                     .readdata
		.coe_exe_start               (leap_profiling_signals_start),                        //    profiling_signals.export
		.coe_exe_end                 (leap_profiling_signals_end),                          //                     .export
		.coe_debug_select            (leap_debug_port_select),                              //           debug_port.export
		.coe_debug_lights            (leap_debug_port_lights)                               //                     .export
	);

	leap_sim_controller #(
		.STARTING_PC (1073741856),
		.N2          (8)
	) leap_sim_control (
		.clk                           (clk_clk),                                                   //         clock.clk
		.reset                         (rst_controller_reset_out_reset),                            //         reset.reset
		.avs_bridge_slave_address      (mm_interconnect_1_leap_sim_control_bridge_slave_address),   //  bridge_slave.address
		.avs_bridge_slave_read         (mm_interconnect_1_leap_sim_control_bridge_slave_read),      //              .read
		.avs_bridge_slave_write        (mm_interconnect_1_leap_sim_control_bridge_slave_write),     //              .write
		.avs_bridge_slave_writedata    (mm_interconnect_1_leap_sim_control_bridge_slave_writedata), //              .writedata
		.avs_bridge_slave_readdata     (mm_interconnect_1_leap_sim_control_bridge_slave_readdata),  //              .readdata
		.avm_bridge_master_readdata    (leap_sim_control_bridge_master_readdata),                   // bridge_master.readdata
		.avm_bridge_master_waitrequest (leap_sim_control_bridge_master_waitrequest),                //              .waitrequest
		.avm_bridge_master_address     (leap_sim_control_bridge_master_address),                    //              .address
		.avm_bridge_master_byteenable  (leap_sim_control_bridge_master_byteenable),                 //              .byteenable
		.avm_bridge_master_read        (leap_sim_control_bridge_master_read),                       //              .read
		.avm_bridge_master_write       (leap_sim_control_bridge_master_write),                      //              .write
		.avm_bridge_master_writedata   (leap_sim_control_bridge_master_writedata)                   //              .writedata
	);

	legup_system_SDRAM sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_1_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_1_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_1_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_1_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_1_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_1_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_1_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_1_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_1_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	tiger_icache_av_1port tiger_icache (
		.clk                                  (clk_clk),                                                   //         clock.clk
		.reset_n                              (~rst_controller_reset_out_reset),                           //         reset.reset_n
		.avs_icache_slave_address             (mm_interconnect_3_tiger_icache_icache_slave_address),       //  icache_slave.address
		.avs_icache_slave_read                (mm_interconnect_3_tiger_icache_icache_slave_read),          //              .read
		.avs_icache_slave_readdata            (mm_interconnect_3_tiger_icache_icache_slave_readdata),      //              .readdata
		.avs_icache_slave_readdatavalid       (mm_interconnect_3_tiger_icache_icache_slave_readdatavalid), //              .readdatavalid
		.avs_icache_slave_waitrequest         (mm_interconnect_3_tiger_icache_icache_slave_waitrequest),   //              .waitrequest
		.avm_icache_master_readdata           (tiger_icache_icache_master_readdata),                       // icache_master.readdata
		.avm_icache_master_readdatavalid      (tiger_icache_icache_master_readdatavalid),                  //              .readdatavalid
		.avm_icache_master_waitrequest        (tiger_icache_icache_master_waitrequest),                    //              .waitrequest
		.avm_icache_master_address            (tiger_icache_icache_master_address),                        //              .address
		.avm_icache_master_beginbursttransfer (tiger_icache_icache_master_beginbursttransfer),             //              .beginbursttransfer
		.avm_icache_master_burstcount         (tiger_icache_icache_master_burstcount),                     //              .burstcount
		.avm_icache_master_read               (tiger_icache_icache_master_read)                            //              .read
	);

	tiger_top #(
		.RESET_ADDRESS (1073741824)
	) tiger_mips (
		.clk                           (clk_clk),                                     //              clock.clk
		.reset                         (rst_controller_001_reset_out_reset),          //              reset.reset
		.avm_instrMaster_address       (tiger_mips_instruction_master_address),       // instruction_master.address
		.avm_instrMaster_read          (tiger_mips_instruction_master_read),          //                   .read
		.avm_instrMaster_write         (tiger_mips_instruction_master_write),         //                   .write
		.avm_instrMaster_writedata     (tiger_mips_instruction_master_writedata),     //                   .writedata
		.avm_instrMaster_byteenable    (tiger_mips_instruction_master_byteenable),    //                   .byteenable
		.avm_instrMaster_readdata      (tiger_mips_instruction_master_readdata),      //                   .readdata
		.avm_instrMaster_waitrequest   (tiger_mips_instruction_master_waitrequest),   //                   .waitrequest
		.avm_instrMaster_readdatavalid (tiger_mips_instruction_master_readdatavalid), //                   .readdatavalid
		.avm_dataMaster_address        (tiger_mips_data_master_address),              //        data_master.address
		.avm_dataMaster_read           (tiger_mips_data_master_read),                 //                   .read
		.avm_dataMaster_write          (tiger_mips_data_master_write),                //                   .write
		.avm_dataMaster_writedata      (tiger_mips_data_master_writedata),            //                   .writedata
		.avm_dataMaster_byteenable     (tiger_mips_data_master_byteenable),           //                   .byteenable
		.avm_dataMaster_readdata       (tiger_mips_data_master_readdata),             //                   .readdata
		.avm_dataMaster_waitrequest    (tiger_mips_data_master_waitrequest),          //                   .waitrequest
		.avm_dataMaster_readdatavalid  (tiger_mips_data_master_readdatavalid)         //                   .readdatavalid
	);

	legup_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                        (clk_clk),                                             //                                      clk_clk.clk
		.Leap_Sim_Control_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                      // Leap_Sim_Control_reset_reset_bridge_in_reset.reset
		.Leap_Sim_Control_bridge_master_address             (leap_sim_control_bridge_master_address),              //               Leap_Sim_Control_bridge_master.address
		.Leap_Sim_Control_bridge_master_waitrequest         (leap_sim_control_bridge_master_waitrequest),          //                                             .waitrequest
		.Leap_Sim_Control_bridge_master_byteenable          (leap_sim_control_bridge_master_byteenable),           //                                             .byteenable
		.Leap_Sim_Control_bridge_master_read                (leap_sim_control_bridge_master_read),                 //                                             .read
		.Leap_Sim_Control_bridge_master_readdata            (leap_sim_control_bridge_master_readdata),             //                                             .readdata
		.Leap_Sim_Control_bridge_master_write               (leap_sim_control_bridge_master_write),                //                                             .write
		.Leap_Sim_Control_bridge_master_writedata           (leap_sim_control_bridge_master_writedata),            //                                             .writedata
		.Leap_Profiler_leapslave_address                    (mm_interconnect_0_leap_profiler_leapslave_address),   //                      Leap_Profiler_leapslave.address
		.Leap_Profiler_leapslave_write                      (mm_interconnect_0_leap_profiler_leapslave_write),     //                                             .write
		.Leap_Profiler_leapslave_read                       (mm_interconnect_0_leap_profiler_leapslave_read),      //                                             .read
		.Leap_Profiler_leapslave_readdata                   (mm_interconnect_0_leap_profiler_leapslave_readdata),  //                                             .readdata
		.Leap_Profiler_leapslave_writedata                  (mm_interconnect_0_leap_profiler_leapslave_writedata)  //                                             .writedata
	);

	legup_system_mm_interconnect_1 mm_interconnect_1 (
		.clk_clk_clk                                               (clk_clk),                                                   //                                             clk_clk.clk
		.DCache_reset_reset_bridge_in_reset_reset                  (rst_controller_reset_out_reset),                            //                  DCache_reset_reset_bridge_in_reset.reset
		.JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset.reset
		.Tiger_MIPS_reset_reset_bridge_in_reset_reset              (rst_controller_001_reset_out_reset),                        //              Tiger_MIPS_reset_reset_bridge_in_reset.reset
		.DCache_cache_master_address                               (dcache_cache_master_address),                               //                                 DCache_cache_master.address
		.DCache_cache_master_waitrequest                           (dcache_cache_master_waitrequest),                           //                                                    .waitrequest
		.DCache_cache_master_burstcount                            (dcache_cache_master_burstcount),                            //                                                    .burstcount
		.DCache_cache_master_byteenable                            (dcache_cache_master_byteenable),                            //                                                    .byteenable
		.DCache_cache_master_read                                  (dcache_cache_master_read),                                  //                                                    .read
		.DCache_cache_master_readdata                              (dcache_cache_master_readdata),                              //                                                    .readdata
		.DCache_cache_master_readdatavalid                         (dcache_cache_master_readdatavalid),                         //                                                    .readdatavalid
		.DCache_cache_master_write                                 (dcache_cache_master_write),                                 //                                                    .write
		.DCache_cache_master_writedata                             (dcache_cache_master_writedata),                             //                                                    .writedata
		.JTAG_to_FPGA_Bridge_master_address                        (jtag_to_fpga_bridge_master_address),                        //                          JTAG_to_FPGA_Bridge_master.address
		.JTAG_to_FPGA_Bridge_master_waitrequest                    (jtag_to_fpga_bridge_master_waitrequest),                    //                                                    .waitrequest
		.JTAG_to_FPGA_Bridge_master_byteenable                     (jtag_to_fpga_bridge_master_byteenable),                     //                                                    .byteenable
		.JTAG_to_FPGA_Bridge_master_read                           (jtag_to_fpga_bridge_master_read),                           //                                                    .read
		.JTAG_to_FPGA_Bridge_master_readdata                       (jtag_to_fpga_bridge_master_readdata),                       //                                                    .readdata
		.JTAG_to_FPGA_Bridge_master_readdatavalid                  (jtag_to_fpga_bridge_master_readdatavalid),                  //                                                    .readdatavalid
		.JTAG_to_FPGA_Bridge_master_write                          (jtag_to_fpga_bridge_master_write),                          //                                                    .write
		.JTAG_to_FPGA_Bridge_master_writedata                      (jtag_to_fpga_bridge_master_writedata),                      //                                                    .writedata
		.Tiger_ICache_icache_master_address                        (tiger_icache_icache_master_address),                        //                          Tiger_ICache_icache_master.address
		.Tiger_ICache_icache_master_waitrequest                    (tiger_icache_icache_master_waitrequest),                    //                                                    .waitrequest
		.Tiger_ICache_icache_master_burstcount                     (tiger_icache_icache_master_burstcount),                     //                                                    .burstcount
		.Tiger_ICache_icache_master_beginbursttransfer             (tiger_icache_icache_master_beginbursttransfer),             //                                                    .beginbursttransfer
		.Tiger_ICache_icache_master_read                           (tiger_icache_icache_master_read),                           //                                                    .read
		.Tiger_ICache_icache_master_readdata                       (tiger_icache_icache_master_readdata),                       //                                                    .readdata
		.Tiger_ICache_icache_master_readdatavalid                  (tiger_icache_icache_master_readdatavalid),                  //                                                    .readdatavalid
		.Tiger_MIPS_data_master_address                            (tiger_mips_data_master_address),                            //                              Tiger_MIPS_data_master.address
		.Tiger_MIPS_data_master_waitrequest                        (tiger_mips_data_master_waitrequest),                        //                                                    .waitrequest
		.Tiger_MIPS_data_master_byteenable                         (tiger_mips_data_master_byteenable),                         //                                                    .byteenable
		.Tiger_MIPS_data_master_read                               (tiger_mips_data_master_read),                               //                                                    .read
		.Tiger_MIPS_data_master_readdata                           (tiger_mips_data_master_readdata),                           //                                                    .readdata
		.Tiger_MIPS_data_master_readdatavalid                      (tiger_mips_data_master_readdatavalid),                      //                                                    .readdatavalid
		.Tiger_MIPS_data_master_write                              (tiger_mips_data_master_write),                              //                                                    .write
		.Tiger_MIPS_data_master_writedata                          (tiger_mips_data_master_writedata),                          //                                                    .writedata
		.DCache_cache_slave_address                                (mm_interconnect_1_dcache_cache_slave_address),              //                                  DCache_cache_slave.address
		.DCache_cache_slave_write                                  (mm_interconnect_1_dcache_cache_slave_write),                //                                                    .write
		.DCache_cache_slave_read                                   (mm_interconnect_1_dcache_cache_slave_read),                 //                                                    .read
		.DCache_cache_slave_readdata                               (mm_interconnect_1_dcache_cache_slave_readdata),             //                                                    .readdata
		.DCache_cache_slave_writedata                              (mm_interconnect_1_dcache_cache_slave_writedata),            //                                                    .writedata
		.DCache_cache_slave_byteenable                             (mm_interconnect_1_dcache_cache_slave_byteenable),           //                                                    .byteenable
		.DCache_cache_slave_readdatavalid                          (mm_interconnect_1_dcache_cache_slave_readdatavalid),        //                                                    .readdatavalid
		.DCache_cache_slave_waitrequest                            (mm_interconnect_1_dcache_cache_slave_waitrequest),          //                                                    .waitrequest
		.JTAG_UART_avalon_jtag_slave_address                       (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                         JTAG_UART_avalon_jtag_slave.address
		.JTAG_UART_avalon_jtag_slave_write                         (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),       //                                                    .write
		.JTAG_UART_avalon_jtag_slave_read                          (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),        //                                                    .read
		.JTAG_UART_avalon_jtag_slave_readdata                      (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                                                    .readdata
		.JTAG_UART_avalon_jtag_slave_writedata                     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                                                    .writedata
		.JTAG_UART_avalon_jtag_slave_waitrequest                   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                                                    .waitrequest
		.JTAG_UART_avalon_jtag_slave_chipselect                    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  //                                                    .chipselect
		.Leap_Sim_Control_bridge_slave_address                     (mm_interconnect_1_leap_sim_control_bridge_slave_address),   //                       Leap_Sim_Control_bridge_slave.address
		.Leap_Sim_Control_bridge_slave_write                       (mm_interconnect_1_leap_sim_control_bridge_slave_write),     //                                                    .write
		.Leap_Sim_Control_bridge_slave_read                        (mm_interconnect_1_leap_sim_control_bridge_slave_read),      //                                                    .read
		.Leap_Sim_Control_bridge_slave_readdata                    (mm_interconnect_1_leap_sim_control_bridge_slave_readdata),  //                                                    .readdata
		.Leap_Sim_Control_bridge_slave_writedata                   (mm_interconnect_1_leap_sim_control_bridge_slave_writedata), //                                                    .writedata
		.SDRAM_s1_address                                          (mm_interconnect_1_sdram_s1_address),                        //                                            SDRAM_s1.address
		.SDRAM_s1_write                                            (mm_interconnect_1_sdram_s1_write),                          //                                                    .write
		.SDRAM_s1_read                                             (mm_interconnect_1_sdram_s1_read),                           //                                                    .read
		.SDRAM_s1_readdata                                         (mm_interconnect_1_sdram_s1_readdata),                       //                                                    .readdata
		.SDRAM_s1_writedata                                        (mm_interconnect_1_sdram_s1_writedata),                      //                                                    .writedata
		.SDRAM_s1_byteenable                                       (mm_interconnect_1_sdram_s1_byteenable),                     //                                                    .byteenable
		.SDRAM_s1_readdatavalid                                    (mm_interconnect_1_sdram_s1_readdatavalid),                  //                                                    .readdatavalid
		.SDRAM_s1_waitrequest                                      (mm_interconnect_1_sdram_s1_waitrequest),                    //                                                    .waitrequest
		.SDRAM_s1_chipselect                                       (mm_interconnect_1_sdram_s1_chipselect)                      //                                                    .chipselect
	);

	legup_system_mm_interconnect_3 mm_interconnect_3 (
		.clk_clk_clk                                     (clk_clk),                                                   //                                   clk_clk.clk
		.Leap_Profiler_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // Leap_Profiler_reset_reset_bridge_in_reset.reset
		.Leap_Profiler_to_memory_address                 (leap_profiler_to_memory_address),                           //                   Leap_Profiler_to_memory.address
		.Leap_Profiler_to_memory_waitrequest             (leap_profiler_to_memory_waitrequest),                       //                                          .waitrequest
		.Leap_Profiler_to_memory_byteenable              (leap_profiler_to_memory_byteenable),                        //                                          .byteenable
		.Leap_Profiler_to_memory_read                    (leap_profiler_to_memory_read),                              //                                          .read
		.Leap_Profiler_to_memory_readdata                (leap_profiler_to_memory_readdata),                          //                                          .readdata
		.Leap_Profiler_to_memory_readdatavalid           (leap_profiler_to_memory_readdatavalid),                     //                                          .readdatavalid
		.Leap_Profiler_to_memory_write                   (leap_profiler_to_memory_write),                             //                                          .write
		.Leap_Profiler_to_memory_writedata               (leap_profiler_to_memory_writedata),                         //                                          .writedata
		.Tiger_ICache_icache_slave_address               (mm_interconnect_3_tiger_icache_icache_slave_address),       //                 Tiger_ICache_icache_slave.address
		.Tiger_ICache_icache_slave_read                  (mm_interconnect_3_tiger_icache_icache_slave_read),          //                                          .read
		.Tiger_ICache_icache_slave_readdata              (mm_interconnect_3_tiger_icache_icache_slave_readdata),      //                                          .readdata
		.Tiger_ICache_icache_slave_readdatavalid         (mm_interconnect_3_tiger_icache_icache_slave_readdatavalid), //                                          .readdatavalid
		.Tiger_ICache_icache_slave_waitrequest           (mm_interconnect_3_tiger_icache_icache_slave_waitrequest)    //                                          .waitrequest
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                           // reset_in0.reset
		.reset_in1      (leap_profiler_leap_processor_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                  //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),       // reset_out.reset
		.reset_req      (),                                         // (terminated)
		.reset_req_in0  (1'b0),                                     // (terminated)
		.reset_req_in1  (1'b0),                                     // (terminated)
		.reset_in2      (1'b0),                                     // (terminated)
		.reset_req_in2  (1'b0),                                     // (terminated)
		.reset_in3      (1'b0),                                     // (terminated)
		.reset_req_in3  (1'b0),                                     // (terminated)
		.reset_in4      (1'b0),                                     // (terminated)
		.reset_req_in4  (1'b0),                                     // (terminated)
		.reset_in5      (1'b0),                                     // (terminated)
		.reset_req_in5  (1'b0),                                     // (terminated)
		.reset_in6      (1'b0),                                     // (terminated)
		.reset_req_in6  (1'b0),                                     // (terminated)
		.reset_in7      (1'b0),                                     // (terminated)
		.reset_req_in7  (1'b0),                                     // (terminated)
		.reset_in8      (1'b0),                                     // (terminated)
		.reset_req_in8  (1'b0),                                     // (terminated)
		.reset_in9      (1'b0),                                     // (terminated)
		.reset_req_in9  (1'b0),                                     // (terminated)
		.reset_in10     (1'b0),                                     // (terminated)
		.reset_req_in10 (1'b0),                                     // (terminated)
		.reset_in11     (1'b0),                                     // (terminated)
		.reset_req_in11 (1'b0),                                     // (terminated)
		.reset_in12     (1'b0),                                     // (terminated)
		.reset_req_in12 (1'b0),                                     // (terminated)
		.reset_in13     (1'b0),                                     // (terminated)
		.reset_req_in13 (1'b0),                                     // (terminated)
		.reset_in14     (1'b0),                                     // (terminated)
		.reset_req_in14 (1'b0),                                     // (terminated)
		.reset_in15     (1'b0),                                     // (terminated)
		.reset_req_in15 (1'b0)                                      // (terminated)
	);

endmodule
