// legup_system_tb.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module legup_system_tb (
		input  wire  oct_rzqin  // oct.rzqin
	);

	wire         legup_system_inst_clk_bfm_clk_clk;         // legup_system_inst_clk_bfm:clk -> [legup_system_inst:clk_clk, legup_system_inst_reset_bfm:clk]
	wire   [0:0] legup_system_inst_ddr3_memory_mem_cas_n;   // legup_system_inst:ddr3_memory_mem_cas_n -> DDR3_SDRAM_mem_model:mem_cas_n
	wire         legup_system_inst_ddr3_memory_mem_reset_n; // legup_system_inst:ddr3_memory_mem_reset_n -> DDR3_SDRAM_mem_model:mem_reset_n
	wire   [2:0] legup_system_inst_ddr3_memory_mem_ba;      // legup_system_inst:ddr3_memory_mem_ba -> DDR3_SDRAM_mem_model:mem_ba
	wire   [0:0] legup_system_inst_ddr3_memory_mem_we_n;    // legup_system_inst:ddr3_memory_mem_we_n -> DDR3_SDRAM_mem_model:mem_we_n
	wire   [0:0] legup_system_inst_ddr3_memory_mem_ck;      // legup_system_inst:ddr3_memory_mem_ck -> DDR3_SDRAM_mem_model:mem_ck
	wire   [7:0] legup_system_inst_ddr3_memory_mem_dm;      // legup_system_inst:ddr3_memory_mem_dm -> DDR3_SDRAM_mem_model:mem_dm
	wire   [7:0] ddr3_sdram_mem_model_memory_mem_dqs;       // [] -> [DDR3_SDRAM_mem_model:mem_dqs, legup_system_inst:ddr3_memory_mem_dqs]
	wire  [63:0] ddr3_sdram_mem_model_memory_mem_dq;        // [] -> [DDR3_SDRAM_mem_model:mem_dq, legup_system_inst:ddr3_memory_mem_dq]
	wire   [0:0] legup_system_inst_ddr3_memory_mem_cs_n;    // legup_system_inst:ddr3_memory_mem_cs_n -> DDR3_SDRAM_mem_model:mem_cs_n
	wire  [13:0] legup_system_inst_ddr3_memory_mem_a;       // legup_system_inst:ddr3_memory_mem_a -> DDR3_SDRAM_mem_model:mem_a
	wire   [0:0] legup_system_inst_ddr3_memory_mem_ras_n;   // legup_system_inst:ddr3_memory_mem_ras_n -> DDR3_SDRAM_mem_model:mem_ras_n
	wire   [7:0] ddr3_sdram_mem_model_memory_mem_dqs_n;     // [] -> [DDR3_SDRAM_mem_model:mem_dqs_n, legup_system_inst:ddr3_memory_mem_dqs_n]
	wire   [0:0] legup_system_inst_ddr3_memory_mem_odt;     // legup_system_inst:ddr3_memory_mem_odt -> DDR3_SDRAM_mem_model:mem_odt
	wire   [0:0] legup_system_inst_ddr3_memory_mem_ck_n;    // legup_system_inst:ddr3_memory_mem_ck_n -> DDR3_SDRAM_mem_model:mem_ck_n
	wire   [0:0] legup_system_inst_ddr3_memory_mem_cke;     // legup_system_inst:ddr3_memory_mem_cke -> DDR3_SDRAM_mem_model:mem_cke
	wire         legup_system_inst_reset_bfm_reset_reset;   // legup_system_inst_reset_bfm:reset -> legup_system_inst:reset_reset_n

	alt_mem_if_ddr3_mem_model_top_ddr3_mem_if_dm_pins_en_mem_if_dqsn_en_udimm #(
		.MEM_IF_ADDR_WIDTH            (14),
		.MEM_IF_ROW_ADDR_WIDTH        (14),
		.MEM_IF_COL_ADDR_WIDTH        (10),
		.MEM_IF_CONTROL_WIDTH         (1),
		.MEM_IF_DQS_WIDTH             (8),
		.MEM_IF_CS_WIDTH              (1),
		.MEM_IF_BANKADDR_WIDTH        (3),
		.MEM_IF_DQ_WIDTH              (64),
		.MEM_IF_CK_WIDTH              (1),
		.MEM_IF_CLK_EN_WIDTH          (1),
		.MEM_TRCD                     (11),
		.MEM_TRTP                     (6),
		.MEM_DQS_TO_CLK_CAPTURE_DELAY (100),
		.MEM_CLK_TO_DQS_CAPTURE_DELAY (100000),
		.MEM_IF_ODT_WIDTH             (1),
		.MEM_IF_LRDIMM_RM             (0),
		.MEM_MIRROR_ADDRESSING_DEC    (0),
		.MEM_REGDIMM_ENABLED          (0),
		.MEM_LRDIMM_ENABLED           (0),
		.DEVICE_DEPTH                 (1),
		.MEM_NUMBER_OF_DIMMS          (1),
		.MEM_NUMBER_OF_RANKS_PER_DIMM (1),
		.MEM_GUARANTEED_WRITE_INIT    (0),
		.MEM_VERBOSE                  (1),
		.REFRESH_BURST_VALIDATION     (0),
		.AP_MODE_EN                   (2'b00),
		.MEM_INIT_EN                  (0),
		.MEM_INIT_FILE                (""),
		.DAT_DATA_WIDTH               (32)
	) ddr3_sdram_mem_model (
		.mem_a       (legup_system_inst_ddr3_memory_mem_a),       // memory.mem_a
		.mem_ba      (legup_system_inst_ddr3_memory_mem_ba),      //       .mem_ba
		.mem_ck      (legup_system_inst_ddr3_memory_mem_ck),      //       .mem_ck
		.mem_ck_n    (legup_system_inst_ddr3_memory_mem_ck_n),    //       .mem_ck_n
		.mem_cke     (legup_system_inst_ddr3_memory_mem_cke),     //       .mem_cke
		.mem_cs_n    (legup_system_inst_ddr3_memory_mem_cs_n),    //       .mem_cs_n
		.mem_dm      (legup_system_inst_ddr3_memory_mem_dm),      //       .mem_dm
		.mem_ras_n   (legup_system_inst_ddr3_memory_mem_ras_n),   //       .mem_ras_n
		.mem_cas_n   (legup_system_inst_ddr3_memory_mem_cas_n),   //       .mem_cas_n
		.mem_we_n    (legup_system_inst_ddr3_memory_mem_we_n),    //       .mem_we_n
		.mem_reset_n (legup_system_inst_ddr3_memory_mem_reset_n), //       .mem_reset_n
		.mem_dq      (ddr3_sdram_mem_model_memory_mem_dq),        //       .mem_dq
		.mem_dqs     (ddr3_sdram_mem_model_memory_mem_dqs),       //       .mem_dqs
		.mem_dqs_n   (ddr3_sdram_mem_model_memory_mem_dqs_n),     //       .mem_dqs_n
		.mem_odt     (legup_system_inst_ddr3_memory_mem_odt)      //       .mem_odt
	);

	legup_system legup_system_inst (
		.clk_clk                       (legup_system_inst_clk_bfm_clk_clk),         //                    clk.clk
		.ddr3_memory_mem_a             (legup_system_inst_ddr3_memory_mem_a),       //            ddr3_memory.mem_a
		.ddr3_memory_mem_ba            (legup_system_inst_ddr3_memory_mem_ba),      //                       .mem_ba
		.ddr3_memory_mem_ck            (legup_system_inst_ddr3_memory_mem_ck),      //                       .mem_ck
		.ddr3_memory_mem_ck_n          (legup_system_inst_ddr3_memory_mem_ck_n),    //                       .mem_ck_n
		.ddr3_memory_mem_cke           (legup_system_inst_ddr3_memory_mem_cke),     //                       .mem_cke
		.ddr3_memory_mem_cs_n          (legup_system_inst_ddr3_memory_mem_cs_n),    //                       .mem_cs_n
		.ddr3_memory_mem_dm            (legup_system_inst_ddr3_memory_mem_dm),      //                       .mem_dm
		.ddr3_memory_mem_ras_n         (legup_system_inst_ddr3_memory_mem_ras_n),   //                       .mem_ras_n
		.ddr3_memory_mem_cas_n         (legup_system_inst_ddr3_memory_mem_cas_n),   //                       .mem_cas_n
		.ddr3_memory_mem_we_n          (legup_system_inst_ddr3_memory_mem_we_n),    //                       .mem_we_n
		.ddr3_memory_mem_reset_n       (legup_system_inst_ddr3_memory_mem_reset_n), //                       .mem_reset_n
		.ddr3_memory_mem_dq            (ddr3_sdram_mem_model_memory_mem_dq),        //                       .mem_dq
		.ddr3_memory_mem_dqs           (ddr3_sdram_mem_model_memory_mem_dqs),       //                       .mem_dqs
		.ddr3_memory_mem_dqs_n         (ddr3_sdram_mem_model_memory_mem_dqs_n),     //                       .mem_dqs_n
		.ddr3_memory_mem_odt           (legup_system_inst_ddr3_memory_mem_odt),     //                       .mem_odt
		.ddr3_oct_rzqin                (oct_rzqin),                                 //               ddr3_oct.rzqin
		.ddr3_status_local_init_done   (),                                          //            ddr3_status.local_init_done
		.ddr3_status_local_cal_success (),                                          //                       .local_cal_success
		.ddr3_status_local_cal_fail    (),                                          //                       .local_cal_fail
		.leap_debug_port_select        (),                                          //        leap_debug_port.select
		.leap_debug_port_lights        (),                                          //                       .lights
		.leap_profiling_signals_start  (),                                          // leap_profiling_signals.start
		.leap_profiling_signals_end    (),                                          //                       .end
		.reset_reset_n                 (legup_system_inst_reset_bfm_reset_reset),   //                  reset.reset_n
		.uart_wire_rxd                 (),                                          //              uart_wire.rxd
		.uart_wire_txd                 ()                                           //                       .txd
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) legup_system_inst_clk_bfm (
		.clk (legup_system_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) legup_system_inst_reset_bfm (
		.reset (legup_system_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (legup_system_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
