module testbench ();

/*****************************************************************************
 *                           Parameter Declarations                          *
 *****************************************************************************/

parameter CLOCK_PERIOD 		= 20;

/*****************************************************************************
 *                             Port Declarations                             *
 *****************************************************************************/
// Inputs

// Bidirectionals

// Outputs

/*****************************************************************************
 *                 Internal Wires and Registers Declarations                 *
 *****************************************************************************/

// Internal Wires

// Internal Registers
reg					clk;
reg					reset;

// State Machine Registers

/*****************************************************************************
 *                         Finite State Machine(s)                           *
 *****************************************************************************/


/*****************************************************************************
 *                             Sequential Logic                              *
 *****************************************************************************/

initial
begin
	clk				<= 1'b0;
end

always
begin : Clock_Generator
	#((CLOCK_PERIOD) / 2) clk = ~clk;
end

initial begin
		reset <= 1'b1;
	#50	reset <= 1'b0;
end

/*****************************************************************************
 *                            Combinational Logic                            *
 *****************************************************************************/


/*****************************************************************************
 *                              Internal Modules                             *
 *****************************************************************************/

sobel sobel (
	// Inputs
	.clk					(clk),
	.reset				(reset),

	.errors				(),
	.done					(),


	.output_mem_data	()
);

endmodule

