// legup_system.v

// Generated using ACDS version 13.0sp1 232 at 2015.05.08.18:58:30

`timescale 1 ps / 1 ps
module legup_system (
		input  wire        clk_clk,                      //                    clk.clk
		input  wire        reset_reset_n,                //                  reset.reset_n
		output wire        leap_profiling_signals_start, // leap_profiling_signals.start
		output wire        leap_profiling_signals_end,   //                       .end
		input  wire [2:0]  leap_debug_port_select,       //        leap_debug_port.select
		output wire [17:0] leap_debug_port_lights,       //                       .lights
		output wire [11:0] sdram_wire_addr,              //             sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                //                       .ba
		output wire        sdram_wire_cas_n,             //                       .cas_n
		output wire        sdram_wire_cke,               //                       .cke
		output wire        sdram_wire_cs_n,              //                       .cs_n
		inout  wire [15:0] sdram_wire_dq,                //                       .dq
		output wire [1:0]  sdram_wire_dqm,               //                       .dqm
		output wire        sdram_wire_ras_n,             //                       .ras_n
		output wire        sdram_wire_we_n,              //                       .we_n
		input  wire        uart_wire_rxd,                //              uart_wire.rxd
		output wire        uart_wire_txd                 //                       .txd
	);

	wire          tiger_mips_instruction_master_waitrequest;                                                          // Leap_Profiler:avs_from_cpu_waitrequest -> Tiger_MIPS:avm_instrMaster_waitrequest
	wire   [31:0] tiger_mips_instruction_master_writedata;                                                            // Tiger_MIPS:avm_instrMaster_writedata -> Leap_Profiler:avs_from_cpu_writedata
	wire   [31:0] tiger_mips_instruction_master_address;                                                              // Tiger_MIPS:avm_instrMaster_address -> Leap_Profiler:avs_from_cpu_address
	wire          tiger_mips_instruction_master_write;                                                                // Tiger_MIPS:avm_instrMaster_write -> Leap_Profiler:avs_from_cpu_write
	wire          tiger_mips_instruction_master_read;                                                                 // Tiger_MIPS:avm_instrMaster_read -> Leap_Profiler:avs_from_cpu_read
	wire   [31:0] tiger_mips_instruction_master_readdata;                                                             // Leap_Profiler:avs_from_cpu_readdata -> Tiger_MIPS:avm_instrMaster_readdata
	wire          tiger_mips_instruction_master_readdatavalid;                                                        // Leap_Profiler:avs_from_cpu_readdatavalid -> Tiger_MIPS:avm_instrMaster_readdatavalid
	wire    [3:0] tiger_mips_instruction_master_byteenable;                                                           // Tiger_MIPS:avm_instrMaster_byteenable -> Leap_Profiler:avs_from_cpu_byteenable
	wire          leap_sim_control_bridge_master_waitrequest;                                                         // Leap_Sim_Control_bridge_master_translator:av_waitrequest -> Leap_Sim_Control:avm_bridge_master_waitrequest
	wire   [31:0] leap_sim_control_bridge_master_writedata;                                                           // Leap_Sim_Control:avm_bridge_master_writedata -> Leap_Sim_Control_bridge_master_translator:av_writedata
	wire   [31:0] leap_sim_control_bridge_master_address;                                                             // Leap_Sim_Control:avm_bridge_master_address -> Leap_Sim_Control_bridge_master_translator:av_address
	wire          leap_sim_control_bridge_master_write;                                                               // Leap_Sim_Control:avm_bridge_master_write -> Leap_Sim_Control_bridge_master_translator:av_write
	wire          leap_sim_control_bridge_master_read;                                                                // Leap_Sim_Control:avm_bridge_master_read -> Leap_Sim_Control_bridge_master_translator:av_read
	wire   [31:0] leap_sim_control_bridge_master_readdata;                                                            // Leap_Sim_Control_bridge_master_translator:av_readdata -> Leap_Sim_Control:avm_bridge_master_readdata
	wire    [3:0] leap_sim_control_bridge_master_byteenable;                                                          // Leap_Sim_Control:avm_bridge_master_byteenable -> Leap_Sim_Control_bridge_master_translator:av_byteenable
	wire          leap_sim_control_bridge_master_translator_avalon_universal_master_0_waitrequest;                    // Leap_Profiler_leapslave_translator:uav_waitrequest -> Leap_Sim_Control_bridge_master_translator:uav_waitrequest
	wire    [2:0] leap_sim_control_bridge_master_translator_avalon_universal_master_0_burstcount;                     // Leap_Sim_Control_bridge_master_translator:uav_burstcount -> Leap_Profiler_leapslave_translator:uav_burstcount
	wire   [31:0] leap_sim_control_bridge_master_translator_avalon_universal_master_0_writedata;                      // Leap_Sim_Control_bridge_master_translator:uav_writedata -> Leap_Profiler_leapslave_translator:uav_writedata
	wire   [31:0] leap_sim_control_bridge_master_translator_avalon_universal_master_0_address;                        // Leap_Sim_Control_bridge_master_translator:uav_address -> Leap_Profiler_leapslave_translator:uav_address
	wire          leap_sim_control_bridge_master_translator_avalon_universal_master_0_lock;                           // Leap_Sim_Control_bridge_master_translator:uav_lock -> Leap_Profiler_leapslave_translator:uav_lock
	wire          leap_sim_control_bridge_master_translator_avalon_universal_master_0_write;                          // Leap_Sim_Control_bridge_master_translator:uav_write -> Leap_Profiler_leapslave_translator:uav_write
	wire          leap_sim_control_bridge_master_translator_avalon_universal_master_0_read;                           // Leap_Sim_Control_bridge_master_translator:uav_read -> Leap_Profiler_leapslave_translator:uav_read
	wire   [31:0] leap_sim_control_bridge_master_translator_avalon_universal_master_0_readdata;                       // Leap_Profiler_leapslave_translator:uav_readdata -> Leap_Sim_Control_bridge_master_translator:uav_readdata
	wire          leap_sim_control_bridge_master_translator_avalon_universal_master_0_debugaccess;                    // Leap_Sim_Control_bridge_master_translator:uav_debugaccess -> Leap_Profiler_leapslave_translator:uav_debugaccess
	wire    [3:0] leap_sim_control_bridge_master_translator_avalon_universal_master_0_byteenable;                     // Leap_Sim_Control_bridge_master_translator:uav_byteenable -> Leap_Profiler_leapslave_translator:uav_byteenable
	wire          leap_sim_control_bridge_master_translator_avalon_universal_master_0_readdatavalid;                  // Leap_Profiler_leapslave_translator:uav_readdatavalid -> Leap_Sim_Control_bridge_master_translator:uav_readdatavalid
	wire   [31:0] leap_profiler_leapslave_translator_avalon_anti_slave_0_writedata;                                   // Leap_Profiler_leapslave_translator:av_writedata -> Leap_Profiler:avs_leapSlave_writedata
	wire   [29:0] leap_profiler_leapslave_translator_avalon_anti_slave_0_address;                                     // Leap_Profiler_leapslave_translator:av_address -> Leap_Profiler:avs_leapSlave_address
	wire          leap_profiler_leapslave_translator_avalon_anti_slave_0_write;                                       // Leap_Profiler_leapslave_translator:av_write -> Leap_Profiler:avs_leapSlave_write
	wire          leap_profiler_leapslave_translator_avalon_anti_slave_0_read;                                        // Leap_Profiler_leapslave_translator:av_read -> Leap_Profiler:avs_leapSlave_read
	wire   [31:0] leap_profiler_leapslave_translator_avalon_anti_slave_0_readdata;                                    // Leap_Profiler:avs_leapSlave_readdata -> Leap_Profiler_leapslave_translator:av_readdata
	wire          leap_profiler_to_memory_waitrequest;                                                                // Leap_Profiler_to_memory_translator:av_waitrequest -> Leap_Profiler:avs_to_memory_waitrequest
	wire   [31:0] leap_profiler_to_memory_writedata;                                                                  // Leap_Profiler:avs_to_memory_writedata -> Leap_Profiler_to_memory_translator:av_writedata
	wire   [31:0] leap_profiler_to_memory_address;                                                                    // Leap_Profiler:avs_to_memory_address -> Leap_Profiler_to_memory_translator:av_address
	wire          leap_profiler_to_memory_write;                                                                      // Leap_Profiler:avs_to_memory_write -> Leap_Profiler_to_memory_translator:av_write
	wire          leap_profiler_to_memory_read;                                                                       // Leap_Profiler:avs_to_memory_read -> Leap_Profiler_to_memory_translator:av_read
	wire   [31:0] leap_profiler_to_memory_readdata;                                                                   // Leap_Profiler_to_memory_translator:av_readdata -> Leap_Profiler:avs_to_memory_readdata
	wire          leap_profiler_to_memory_readdatavalid;                                                              // Leap_Profiler_to_memory_translator:av_readdatavalid -> Leap_Profiler:avs_to_memory_readdatavalid
	wire    [3:0] leap_profiler_to_memory_byteenable;                                                                 // Leap_Profiler:avs_to_memory_byteenable -> Leap_Profiler_to_memory_translator:av_byteenable
	wire          leap_profiler_to_memory_translator_avalon_universal_master_0_waitrequest;                           // Tiger_ICache_icache_slave_translator:uav_waitrequest -> Leap_Profiler_to_memory_translator:uav_waitrequest
	wire    [2:0] leap_profiler_to_memory_translator_avalon_universal_master_0_burstcount;                            // Leap_Profiler_to_memory_translator:uav_burstcount -> Tiger_ICache_icache_slave_translator:uav_burstcount
	wire   [31:0] leap_profiler_to_memory_translator_avalon_universal_master_0_writedata;                             // Leap_Profiler_to_memory_translator:uav_writedata -> Tiger_ICache_icache_slave_translator:uav_writedata
	wire   [31:0] leap_profiler_to_memory_translator_avalon_universal_master_0_address;                               // Leap_Profiler_to_memory_translator:uav_address -> Tiger_ICache_icache_slave_translator:uav_address
	wire          leap_profiler_to_memory_translator_avalon_universal_master_0_lock;                                  // Leap_Profiler_to_memory_translator:uav_lock -> Tiger_ICache_icache_slave_translator:uav_lock
	wire          leap_profiler_to_memory_translator_avalon_universal_master_0_write;                                 // Leap_Profiler_to_memory_translator:uav_write -> Tiger_ICache_icache_slave_translator:uav_write
	wire          leap_profiler_to_memory_translator_avalon_universal_master_0_read;                                  // Leap_Profiler_to_memory_translator:uav_read -> Tiger_ICache_icache_slave_translator:uav_read
	wire   [31:0] leap_profiler_to_memory_translator_avalon_universal_master_0_readdata;                              // Tiger_ICache_icache_slave_translator:uav_readdata -> Leap_Profiler_to_memory_translator:uav_readdata
	wire          leap_profiler_to_memory_translator_avalon_universal_master_0_debugaccess;                           // Leap_Profiler_to_memory_translator:uav_debugaccess -> Tiger_ICache_icache_slave_translator:uav_debugaccess
	wire    [3:0] leap_profiler_to_memory_translator_avalon_universal_master_0_byteenable;                            // Leap_Profiler_to_memory_translator:uav_byteenable -> Tiger_ICache_icache_slave_translator:uav_byteenable
	wire          leap_profiler_to_memory_translator_avalon_universal_master_0_readdatavalid;                         // Tiger_ICache_icache_slave_translator:uav_readdatavalid -> Leap_Profiler_to_memory_translator:uav_readdatavalid
	wire          tiger_icache_icache_slave_translator_avalon_anti_slave_0_waitrequest;                               // Tiger_ICache:avs_icache_slave_waitrequest -> Tiger_ICache_icache_slave_translator:av_waitrequest
	wire   [29:0] tiger_icache_icache_slave_translator_avalon_anti_slave_0_address;                                   // Tiger_ICache_icache_slave_translator:av_address -> Tiger_ICache:avs_icache_slave_address
	wire          tiger_icache_icache_slave_translator_avalon_anti_slave_0_read;                                      // Tiger_ICache_icache_slave_translator:av_read -> Tiger_ICache:avs_icache_slave_read
	wire   [31:0] tiger_icache_icache_slave_translator_avalon_anti_slave_0_readdata;                                  // Tiger_ICache:avs_icache_slave_readdata -> Tiger_ICache_icache_slave_translator:av_readdata
	wire          tiger_icache_icache_slave_translator_avalon_anti_slave_0_readdatavalid;                             // Tiger_ICache:avs_icache_slave_readdatavalid -> Tiger_ICache_icache_slave_translator:av_readdatavalid
	wire          tiger_mips_data_master_waitrequest;                                                                 // Tiger_MIPS_data_master_translator:av_waitrequest -> Tiger_MIPS:avm_dataMaster_waitrequest
	wire   [31:0] tiger_mips_data_master_writedata;                                                                   // Tiger_MIPS:avm_dataMaster_writedata -> Tiger_MIPS_data_master_translator:av_writedata
	wire   [31:0] tiger_mips_data_master_address;                                                                     // Tiger_MIPS:avm_dataMaster_address -> Tiger_MIPS_data_master_translator:av_address
	wire          tiger_mips_data_master_write;                                                                       // Tiger_MIPS:avm_dataMaster_write -> Tiger_MIPS_data_master_translator:av_write
	wire          tiger_mips_data_master_read;                                                                        // Tiger_MIPS:avm_dataMaster_read -> Tiger_MIPS_data_master_translator:av_read
	wire   [31:0] tiger_mips_data_master_readdata;                                                                    // Tiger_MIPS_data_master_translator:av_readdata -> Tiger_MIPS:avm_dataMaster_readdata
	wire          tiger_mips_data_master_readdatavalid;                                                               // Tiger_MIPS_data_master_translator:av_readdatavalid -> Tiger_MIPS:avm_dataMaster_readdatavalid
	wire    [3:0] tiger_mips_data_master_byteenable;                                                                  // Tiger_MIPS:avm_dataMaster_byteenable -> Tiger_MIPS_data_master_translator:av_byteenable
	wire          jtag_to_fpga_bridge_master_waitrequest;                                                             // JTAG_to_FPGA_Bridge_master_translator:av_waitrequest -> JTAG_to_FPGA_Bridge:master_waitrequest
	wire   [31:0] jtag_to_fpga_bridge_master_writedata;                                                               // JTAG_to_FPGA_Bridge:master_writedata -> JTAG_to_FPGA_Bridge_master_translator:av_writedata
	wire   [31:0] jtag_to_fpga_bridge_master_address;                                                                 // JTAG_to_FPGA_Bridge:master_address -> JTAG_to_FPGA_Bridge_master_translator:av_address
	wire          jtag_to_fpga_bridge_master_write;                                                                   // JTAG_to_FPGA_Bridge:master_write -> JTAG_to_FPGA_Bridge_master_translator:av_write
	wire          jtag_to_fpga_bridge_master_read;                                                                    // JTAG_to_FPGA_Bridge:master_read -> JTAG_to_FPGA_Bridge_master_translator:av_read
	wire   [31:0] jtag_to_fpga_bridge_master_readdata;                                                                // JTAG_to_FPGA_Bridge_master_translator:av_readdata -> JTAG_to_FPGA_Bridge:master_readdata
	wire    [3:0] jtag_to_fpga_bridge_master_byteenable;                                                              // JTAG_to_FPGA_Bridge:master_byteenable -> JTAG_to_FPGA_Bridge_master_translator:av_byteenable
	wire          jtag_to_fpga_bridge_master_readdatavalid;                                                           // JTAG_to_FPGA_Bridge_master_translator:av_readdatavalid -> JTAG_to_FPGA_Bridge:master_readdatavalid
	wire    [5:0] tiger_icache_icache_master_burstcount;                                                              // Tiger_ICache:avm_icache_master_burstcount -> Tiger_ICache_icache_master_translator:av_burstcount
	wire          tiger_icache_icache_master_waitrequest;                                                             // Tiger_ICache_icache_master_translator:av_waitrequest -> Tiger_ICache:avm_icache_master_waitrequest
	wire   [31:0] tiger_icache_icache_master_address;                                                                 // Tiger_ICache:avm_icache_master_address -> Tiger_ICache_icache_master_translator:av_address
	wire          tiger_icache_icache_master_read;                                                                    // Tiger_ICache:avm_icache_master_read -> Tiger_ICache_icache_master_translator:av_read
	wire          tiger_icache_icache_master_beginbursttransfer;                                                      // Tiger_ICache:avm_icache_master_beginbursttransfer -> Tiger_ICache_icache_master_translator:av_beginbursttransfer
	wire   [31:0] tiger_icache_icache_master_readdata;                                                                // Tiger_ICache_icache_master_translator:av_readdata -> Tiger_ICache:avm_icache_master_readdata
	wire          tiger_icache_icache_master_readdatavalid;                                                           // Tiger_ICache_icache_master_translator:av_readdatavalid -> Tiger_ICache:avm_icache_master_readdatavalid
	wire    [2:0] dcache_cache_master_burstcount;                                                                     // DCache:avm_cache_burstcount -> DCache_cache_master_translator:av_burstcount
	wire          dcache_cache_master_waitrequest;                                                                    // DCache_cache_master_translator:av_waitrequest -> DCache:avm_cache_waitrequest
	wire   [31:0] dcache_cache_master_writedata;                                                                      // DCache:avm_cache_writedata -> DCache_cache_master_translator:av_writedata
	wire   [31:0] dcache_cache_master_address;                                                                        // DCache:avm_cache_address -> DCache_cache_master_translator:av_address
	wire          dcache_cache_master_write;                                                                          // DCache:avm_cache_write -> DCache_cache_master_translator:av_write
	wire          dcache_cache_master_read;                                                                           // DCache:avm_cache_read -> DCache_cache_master_translator:av_read
	wire   [31:0] dcache_cache_master_readdata;                                                                       // DCache_cache_master_translator:av_readdata -> DCache:avm_cache_readdata
	wire    [3:0] dcache_cache_master_byteenable;                                                                     // DCache:avm_cache_byteenable -> DCache_cache_master_translator:av_byteenable
	wire          dcache_cache_master_readdatavalid;                                                                  // DCache_cache_master_translator:av_readdatavalid -> DCache:avm_cache_readdatavalid
	wire          dcache_cache_slave_translator_avalon_anti_slave_0_waitrequest;                                      // DCache:avs_cache_waitrequest -> DCache_cache_slave_translator:av_waitrequest
	wire   [31:0] dcache_cache_slave_translator_avalon_anti_slave_0_writedata;                                        // DCache_cache_slave_translator:av_writedata -> DCache:avs_cache_writedata
	wire   [30:0] dcache_cache_slave_translator_avalon_anti_slave_0_address;                                          // DCache_cache_slave_translator:av_address -> DCache:avs_cache_address
	wire          dcache_cache_slave_translator_avalon_anti_slave_0_write;                                            // DCache_cache_slave_translator:av_write -> DCache:avs_cache_write
	wire          dcache_cache_slave_translator_avalon_anti_slave_0_read;                                             // DCache_cache_slave_translator:av_read -> DCache:avs_cache_read
	wire   [31:0] dcache_cache_slave_translator_avalon_anti_slave_0_readdata;                                         // DCache:avs_cache_readdata -> DCache_cache_slave_translator:av_readdata
	wire          dcache_cache_slave_translator_avalon_anti_slave_0_readdatavalid;                                    // DCache:avs_cache_readdatavalid -> DCache_cache_slave_translator:av_readdatavalid
	wire    [3:0] dcache_cache_slave_translator_avalon_anti_slave_0_byteenable;                                       // DCache_cache_slave_translator:av_byteenable -> DCache:avs_cache_byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                             // JTAG_UART:av_waitrequest -> JTAG_UART_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                               // JTAG_UART_avalon_jtag_slave_translator:av_writedata -> JTAG_UART:av_writedata
	wire    [0:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                 // JTAG_UART_avalon_jtag_slave_translator:av_address -> JTAG_UART:av_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                              // JTAG_UART_avalon_jtag_slave_translator:av_chipselect -> JTAG_UART:av_chipselect
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                   // JTAG_UART_avalon_jtag_slave_translator:av_write -> JTAG_UART:av_write_n
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                    // JTAG_UART_avalon_jtag_slave_translator:av_read -> JTAG_UART:av_read_n
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                // JTAG_UART:av_readdata -> JTAG_UART_avalon_jtag_slave_translator:av_readdata
	wire   [15:0] uart_s1_translator_avalon_anti_slave_0_writedata;                                                   // UART_s1_translator:av_writedata -> UART:writedata
	wire    [2:0] uart_s1_translator_avalon_anti_slave_0_address;                                                     // UART_s1_translator:av_address -> UART:address
	wire          uart_s1_translator_avalon_anti_slave_0_chipselect;                                                  // UART_s1_translator:av_chipselect -> UART:chipselect
	wire          uart_s1_translator_avalon_anti_slave_0_write;                                                       // UART_s1_translator:av_write -> UART:write_n
	wire          uart_s1_translator_avalon_anti_slave_0_read;                                                        // UART_s1_translator:av_read -> UART:read_n
	wire   [15:0] uart_s1_translator_avalon_anti_slave_0_readdata;                                                    // UART:readdata -> UART_s1_translator:av_readdata
	wire          uart_s1_translator_avalon_anti_slave_0_begintransfer;                                               // UART_s1_translator:av_begintransfer -> UART:begintransfer
	wire   [31:0] leap_sim_control_bridge_slave_translator_avalon_anti_slave_0_writedata;                             // Leap_Sim_Control_bridge_slave_translator:av_writedata -> Leap_Sim_Control:avs_bridge_slave_writedata
	wire    [7:0] leap_sim_control_bridge_slave_translator_avalon_anti_slave_0_address;                               // Leap_Sim_Control_bridge_slave_translator:av_address -> Leap_Sim_Control:avs_bridge_slave_address
	wire          leap_sim_control_bridge_slave_translator_avalon_anti_slave_0_write;                                 // Leap_Sim_Control_bridge_slave_translator:av_write -> Leap_Sim_Control:avs_bridge_slave_write
	wire          leap_sim_control_bridge_slave_translator_avalon_anti_slave_0_read;                                  // Leap_Sim_Control_bridge_slave_translator:av_read -> Leap_Sim_Control:avs_bridge_slave_read
	wire   [31:0] leap_sim_control_bridge_slave_translator_avalon_anti_slave_0_readdata;                              // Leap_Sim_Control:avs_bridge_slave_readdata -> Leap_Sim_Control_bridge_slave_translator:av_readdata
	wire          sdram_s1_translator_avalon_anti_slave_0_waitrequest;                                                // SDRAM:za_waitrequest -> SDRAM_s1_translator:av_waitrequest
	wire   [15:0] sdram_s1_translator_avalon_anti_slave_0_writedata;                                                  // SDRAM_s1_translator:av_writedata -> SDRAM:az_data
	wire   [21:0] sdram_s1_translator_avalon_anti_slave_0_address;                                                    // SDRAM_s1_translator:av_address -> SDRAM:az_addr
	wire          sdram_s1_translator_avalon_anti_slave_0_chipselect;                                                 // SDRAM_s1_translator:av_chipselect -> SDRAM:az_cs
	wire          sdram_s1_translator_avalon_anti_slave_0_write;                                                      // SDRAM_s1_translator:av_write -> SDRAM:az_wr_n
	wire          sdram_s1_translator_avalon_anti_slave_0_read;                                                       // SDRAM_s1_translator:av_read -> SDRAM:az_rd_n
	wire   [15:0] sdram_s1_translator_avalon_anti_slave_0_readdata;                                                   // SDRAM:za_data -> SDRAM_s1_translator:av_readdata
	wire          sdram_s1_translator_avalon_anti_slave_0_readdatavalid;                                              // SDRAM:za_valid -> SDRAM_s1_translator:av_readdatavalid
	wire    [1:0] sdram_s1_translator_avalon_anti_slave_0_byteenable;                                                 // SDRAM_s1_translator:av_byteenable -> SDRAM:az_be_n
	wire          tiger_mips_data_master_translator_avalon_universal_master_0_waitrequest;                            // Tiger_MIPS_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> Tiger_MIPS_data_master_translator:uav_waitrequest
	wire    [2:0] tiger_mips_data_master_translator_avalon_universal_master_0_burstcount;                             // Tiger_MIPS_data_master_translator:uav_burstcount -> Tiger_MIPS_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] tiger_mips_data_master_translator_avalon_universal_master_0_writedata;                              // Tiger_MIPS_data_master_translator:uav_writedata -> Tiger_MIPS_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] tiger_mips_data_master_translator_avalon_universal_master_0_address;                                // Tiger_MIPS_data_master_translator:uav_address -> Tiger_MIPS_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          tiger_mips_data_master_translator_avalon_universal_master_0_lock;                                   // Tiger_MIPS_data_master_translator:uav_lock -> Tiger_MIPS_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          tiger_mips_data_master_translator_avalon_universal_master_0_write;                                  // Tiger_MIPS_data_master_translator:uav_write -> Tiger_MIPS_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          tiger_mips_data_master_translator_avalon_universal_master_0_read;                                   // Tiger_MIPS_data_master_translator:uav_read -> Tiger_MIPS_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] tiger_mips_data_master_translator_avalon_universal_master_0_readdata;                               // Tiger_MIPS_data_master_translator_avalon_universal_master_0_agent:av_readdata -> Tiger_MIPS_data_master_translator:uav_readdata
	wire          tiger_mips_data_master_translator_avalon_universal_master_0_debugaccess;                            // Tiger_MIPS_data_master_translator:uav_debugaccess -> Tiger_MIPS_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] tiger_mips_data_master_translator_avalon_universal_master_0_byteenable;                             // Tiger_MIPS_data_master_translator:uav_byteenable -> Tiger_MIPS_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          tiger_mips_data_master_translator_avalon_universal_master_0_readdatavalid;                          // Tiger_MIPS_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> Tiger_MIPS_data_master_translator:uav_readdatavalid
	wire          jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_waitrequest;                        // JTAG_to_FPGA_Bridge_master_translator_avalon_universal_master_0_agent:av_waitrequest -> JTAG_to_FPGA_Bridge_master_translator:uav_waitrequest
	wire    [2:0] jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_burstcount;                         // JTAG_to_FPGA_Bridge_master_translator:uav_burstcount -> JTAG_to_FPGA_Bridge_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_writedata;                          // JTAG_to_FPGA_Bridge_master_translator:uav_writedata -> JTAG_to_FPGA_Bridge_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_address;                            // JTAG_to_FPGA_Bridge_master_translator:uav_address -> JTAG_to_FPGA_Bridge_master_translator_avalon_universal_master_0_agent:av_address
	wire          jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_lock;                               // JTAG_to_FPGA_Bridge_master_translator:uav_lock -> JTAG_to_FPGA_Bridge_master_translator_avalon_universal_master_0_agent:av_lock
	wire          jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_write;                              // JTAG_to_FPGA_Bridge_master_translator:uav_write -> JTAG_to_FPGA_Bridge_master_translator_avalon_universal_master_0_agent:av_write
	wire          jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_read;                               // JTAG_to_FPGA_Bridge_master_translator:uav_read -> JTAG_to_FPGA_Bridge_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_readdata;                           // JTAG_to_FPGA_Bridge_master_translator_avalon_universal_master_0_agent:av_readdata -> JTAG_to_FPGA_Bridge_master_translator:uav_readdata
	wire          jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_debugaccess;                        // JTAG_to_FPGA_Bridge_master_translator:uav_debugaccess -> JTAG_to_FPGA_Bridge_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_byteenable;                         // JTAG_to_FPGA_Bridge_master_translator:uav_byteenable -> JTAG_to_FPGA_Bridge_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_readdatavalid;                      // JTAG_to_FPGA_Bridge_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> JTAG_to_FPGA_Bridge_master_translator:uav_readdatavalid
	wire          tiger_icache_icache_master_translator_avalon_universal_master_0_waitrequest;                        // Tiger_ICache_icache_master_translator_avalon_universal_master_0_agent:av_waitrequest -> Tiger_ICache_icache_master_translator:uav_waitrequest
	wire    [7:0] tiger_icache_icache_master_translator_avalon_universal_master_0_burstcount;                         // Tiger_ICache_icache_master_translator:uav_burstcount -> Tiger_ICache_icache_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] tiger_icache_icache_master_translator_avalon_universal_master_0_writedata;                          // Tiger_ICache_icache_master_translator:uav_writedata -> Tiger_ICache_icache_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] tiger_icache_icache_master_translator_avalon_universal_master_0_address;                            // Tiger_ICache_icache_master_translator:uav_address -> Tiger_ICache_icache_master_translator_avalon_universal_master_0_agent:av_address
	wire          tiger_icache_icache_master_translator_avalon_universal_master_0_lock;                               // Tiger_ICache_icache_master_translator:uav_lock -> Tiger_ICache_icache_master_translator_avalon_universal_master_0_agent:av_lock
	wire          tiger_icache_icache_master_translator_avalon_universal_master_0_write;                              // Tiger_ICache_icache_master_translator:uav_write -> Tiger_ICache_icache_master_translator_avalon_universal_master_0_agent:av_write
	wire          tiger_icache_icache_master_translator_avalon_universal_master_0_read;                               // Tiger_ICache_icache_master_translator:uav_read -> Tiger_ICache_icache_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] tiger_icache_icache_master_translator_avalon_universal_master_0_readdata;                           // Tiger_ICache_icache_master_translator_avalon_universal_master_0_agent:av_readdata -> Tiger_ICache_icache_master_translator:uav_readdata
	wire          tiger_icache_icache_master_translator_avalon_universal_master_0_debugaccess;                        // Tiger_ICache_icache_master_translator:uav_debugaccess -> Tiger_ICache_icache_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] tiger_icache_icache_master_translator_avalon_universal_master_0_byteenable;                         // Tiger_ICache_icache_master_translator:uav_byteenable -> Tiger_ICache_icache_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          tiger_icache_icache_master_translator_avalon_universal_master_0_readdatavalid;                      // Tiger_ICache_icache_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> Tiger_ICache_icache_master_translator:uav_readdatavalid
	wire          dcache_cache_master_translator_avalon_universal_master_0_waitrequest;                               // DCache_cache_master_translator_avalon_universal_master_0_agent:av_waitrequest -> DCache_cache_master_translator:uav_waitrequest
	wire    [4:0] dcache_cache_master_translator_avalon_universal_master_0_burstcount;                                // DCache_cache_master_translator:uav_burstcount -> DCache_cache_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] dcache_cache_master_translator_avalon_universal_master_0_writedata;                                 // DCache_cache_master_translator:uav_writedata -> DCache_cache_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] dcache_cache_master_translator_avalon_universal_master_0_address;                                   // DCache_cache_master_translator:uav_address -> DCache_cache_master_translator_avalon_universal_master_0_agent:av_address
	wire          dcache_cache_master_translator_avalon_universal_master_0_lock;                                      // DCache_cache_master_translator:uav_lock -> DCache_cache_master_translator_avalon_universal_master_0_agent:av_lock
	wire          dcache_cache_master_translator_avalon_universal_master_0_write;                                     // DCache_cache_master_translator:uav_write -> DCache_cache_master_translator_avalon_universal_master_0_agent:av_write
	wire          dcache_cache_master_translator_avalon_universal_master_0_read;                                      // DCache_cache_master_translator:uav_read -> DCache_cache_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] dcache_cache_master_translator_avalon_universal_master_0_readdata;                                  // DCache_cache_master_translator_avalon_universal_master_0_agent:av_readdata -> DCache_cache_master_translator:uav_readdata
	wire          dcache_cache_master_translator_avalon_universal_master_0_debugaccess;                               // DCache_cache_master_translator:uav_debugaccess -> DCache_cache_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] dcache_cache_master_translator_avalon_universal_master_0_byteenable;                                // DCache_cache_master_translator:uav_byteenable -> DCache_cache_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          dcache_cache_master_translator_avalon_universal_master_0_readdatavalid;                             // DCache_cache_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> DCache_cache_master_translator:uav_readdatavalid
	wire          dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // DCache_cache_slave_translator:uav_waitrequest -> DCache_cache_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // DCache_cache_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> DCache_cache_slave_translator:uav_burstcount
	wire   [31:0] dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                          // DCache_cache_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> DCache_cache_slave_translator:uav_writedata
	wire   [31:0] dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_address;                            // DCache_cache_slave_translator_avalon_universal_slave_0_agent:m0_address -> DCache_cache_slave_translator:uav_address
	wire          dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_write;                              // DCache_cache_slave_translator_avalon_universal_slave_0_agent:m0_write -> DCache_cache_slave_translator:uav_write
	wire          dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_lock;                               // DCache_cache_slave_translator_avalon_universal_slave_0_agent:m0_lock -> DCache_cache_slave_translator:uav_lock
	wire          dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_read;                               // DCache_cache_slave_translator_avalon_universal_slave_0_agent:m0_read -> DCache_cache_slave_translator:uav_read
	wire   [31:0] dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                           // DCache_cache_slave_translator:uav_readdata -> DCache_cache_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // DCache_cache_slave_translator:uav_readdatavalid -> DCache_cache_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // DCache_cache_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> DCache_cache_slave_translator:uav_debugaccess
	wire    [3:0] dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // DCache_cache_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> DCache_cache_slave_translator:uav_byteenable
	wire          dcache_cache_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // DCache_cache_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> DCache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          dcache_cache_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // DCache_cache_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> DCache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          dcache_cache_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // DCache_cache_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> DCache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [108:0] dcache_cache_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                        // DCache_cache_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> DCache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          dcache_cache_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // DCache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> DCache_cache_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          dcache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // DCache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> DCache_cache_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          dcache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // DCache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> DCache_cache_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          dcache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // DCache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> DCache_cache_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [108:0] dcache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // DCache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> DCache_cache_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          dcache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // DCache_cache_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> DCache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          dcache_cache_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // DCache_cache_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> DCache_cache_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] dcache_cache_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // DCache_cache_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> DCache_cache_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          dcache_cache_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // DCache_cache_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> DCache_cache_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;               // JTAG_UART_avalon_jtag_slave_translator:uav_waitrequest -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> JTAG_UART_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                 // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> JTAG_UART_avalon_jtag_slave_translator:uav_writedata
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                   // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> JTAG_UART_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                     // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> JTAG_UART_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                      // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> JTAG_UART_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                      // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> JTAG_UART_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                  // JTAG_UART_avalon_jtag_slave_translator:uav_readdata -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;             // JTAG_UART_avalon_jtag_slave_translator:uav_readdatavalid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;               // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> JTAG_UART_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> JTAG_UART_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;        // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;              // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;      // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [108:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;               // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;              // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;     // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;           // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;   // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [108:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;            // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;           // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;         // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;          // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;         // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          uart_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // UART_s1_translator:uav_waitrequest -> UART_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] uart_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // UART_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> UART_s1_translator:uav_burstcount
	wire   [31:0] uart_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // UART_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> UART_s1_translator:uav_writedata
	wire   [31:0] uart_s1_translator_avalon_universal_slave_0_agent_m0_address;                                       // UART_s1_translator_avalon_universal_slave_0_agent:m0_address -> UART_s1_translator:uav_address
	wire          uart_s1_translator_avalon_universal_slave_0_agent_m0_write;                                         // UART_s1_translator_avalon_universal_slave_0_agent:m0_write -> UART_s1_translator:uav_write
	wire          uart_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                          // UART_s1_translator_avalon_universal_slave_0_agent:m0_lock -> UART_s1_translator:uav_lock
	wire          uart_s1_translator_avalon_universal_slave_0_agent_m0_read;                                          // UART_s1_translator_avalon_universal_slave_0_agent:m0_read -> UART_s1_translator:uav_read
	wire   [31:0] uart_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // UART_s1_translator:uav_readdata -> UART_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          uart_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // UART_s1_translator:uav_readdatavalid -> UART_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          uart_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // UART_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> UART_s1_translator:uav_debugaccess
	wire    [3:0] uart_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // UART_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> UART_s1_translator:uav_byteenable
	wire          uart_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // UART_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> UART_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          uart_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // UART_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> UART_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          uart_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // UART_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> UART_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [108:0] uart_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // UART_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> UART_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          uart_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // UART_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> UART_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // UART_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> UART_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // UART_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> UART_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // UART_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> UART_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [108:0] uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // UART_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> UART_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // UART_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> UART_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // UART_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> UART_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // UART_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> UART_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // UART_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> UART_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Leap_Sim_Control_bridge_slave_translator:uav_waitrequest -> Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Leap_Sim_Control_bridge_slave_translator:uav_burstcount
	wire   [31:0] leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Leap_Sim_Control_bridge_slave_translator:uav_writedata
	wire   [31:0] leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:m0_address -> Leap_Sim_Control_bridge_slave_translator:uav_address
	wire          leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:m0_write -> Leap_Sim_Control_bridge_slave_translator:uav_write
	wire          leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Leap_Sim_Control_bridge_slave_translator:uav_lock
	wire          leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:m0_read -> Leap_Sim_Control_bridge_slave_translator:uav_read
	wire   [31:0] leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // Leap_Sim_Control_bridge_slave_translator:uav_readdata -> Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Leap_Sim_Control_bridge_slave_translator:uav_readdatavalid -> Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Leap_Sim_Control_bridge_slave_translator:uav_debugaccess
	wire    [3:0] leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Leap_Sim_Control_bridge_slave_translator:uav_byteenable
	wire          leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [108:0] leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [108:0] leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // SDRAM_s1_translator:uav_waitrequest -> SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> SDRAM_s1_translator:uav_burstcount
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> SDRAM_s1_translator:uav_writedata
	wire   [31:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_address -> SDRAM_s1_translator:uav_address
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_write -> SDRAM_s1_translator:uav_write
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_lock -> SDRAM_s1_translator:uav_lock
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_read -> SDRAM_s1_translator:uav_read
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // SDRAM_s1_translator:uav_readdata -> SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // SDRAM_s1_translator:uav_readdatavalid -> SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SDRAM_s1_translator:uav_debugaccess
	wire    [1:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // SDRAM_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> SDRAM_s1_translator:uav_byteenable
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [90:0] sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [90:0] sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // SDRAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // SDRAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SDRAM_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [17:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // SDRAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SDRAM_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // SDRAM_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                            // SDRAM_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [17:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                             // SDRAM_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                            // SDRAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SDRAM_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          tiger_mips_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                   // Tiger_MIPS_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          tiger_mips_data_master_translator_avalon_universal_master_0_agent_cp_valid;                         // Tiger_MIPS_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          tiger_mips_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                 // Tiger_MIPS_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [107:0] tiger_mips_data_master_translator_avalon_universal_master_0_agent_cp_data;                          // Tiger_MIPS_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          tiger_mips_data_master_translator_avalon_universal_master_0_agent_cp_ready;                         // addr_router:sink_ready -> Tiger_MIPS_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_agent_cp_endofpacket;               // JTAG_to_FPGA_Bridge_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_agent_cp_valid;                     // JTAG_to_FPGA_Bridge_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_agent_cp_startofpacket;             // JTAG_to_FPGA_Bridge_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [107:0] jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_agent_cp_data;                      // JTAG_to_FPGA_Bridge_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_agent_cp_ready;                     // addr_router_001:sink_ready -> JTAG_to_FPGA_Bridge_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          tiger_icache_icache_master_translator_avalon_universal_master_0_agent_cp_endofpacket;               // Tiger_ICache_icache_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          tiger_icache_icache_master_translator_avalon_universal_master_0_agent_cp_valid;                     // Tiger_ICache_icache_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          tiger_icache_icache_master_translator_avalon_universal_master_0_agent_cp_startofpacket;             // Tiger_ICache_icache_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [107:0] tiger_icache_icache_master_translator_avalon_universal_master_0_agent_cp_data;                      // Tiger_ICache_icache_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          tiger_icache_icache_master_translator_avalon_universal_master_0_agent_cp_ready;                     // addr_router_002:sink_ready -> Tiger_ICache_icache_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          dcache_cache_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                      // DCache_cache_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire          dcache_cache_master_translator_avalon_universal_master_0_agent_cp_valid;                            // DCache_cache_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire          dcache_cache_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                    // DCache_cache_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire  [107:0] dcache_cache_master_translator_avalon_universal_master_0_agent_cp_data;                             // DCache_cache_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire          dcache_cache_master_translator_avalon_universal_master_0_agent_cp_ready;                            // addr_router_003:sink_ready -> DCache_cache_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          dcache_cache_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // DCache_cache_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          dcache_cache_slave_translator_avalon_universal_slave_0_agent_rp_valid;                              // DCache_cache_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          dcache_cache_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // DCache_cache_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [107:0] dcache_cache_slave_translator_avalon_universal_slave_0_agent_rp_data;                               // DCache_cache_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          dcache_cache_slave_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router:sink_ready -> DCache_cache_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;               // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                     // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;             // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [107:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                      // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                     // id_router_001:sink_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          uart_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // UART_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          uart_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                         // UART_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          uart_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // UART_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [107:0] uart_s1_translator_avalon_universal_slave_0_agent_rp_data;                                          // UART_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          uart_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_002:sink_ready -> UART_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [107:0] leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_003:sink_ready -> Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // SDRAM_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // SDRAM_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // SDRAM_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire   [89:0] sdram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // SDRAM_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_004:sink_ready -> SDRAM_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_src_endofpacket;                                                                        // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                              // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                                      // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [107:0] addr_router_src_data;                                                                               // addr_router:src_data -> limiter:cmd_sink_data
	wire    [4:0] addr_router_src_channel;                                                                            // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                              // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                        // limiter:rsp_src_endofpacket -> Tiger_MIPS_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                              // limiter:rsp_src_valid -> Tiger_MIPS_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                      // limiter:rsp_src_startofpacket -> Tiger_MIPS_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [107:0] limiter_rsp_src_data;                                                                               // limiter:rsp_src_data -> Tiger_MIPS_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [4:0] limiter_rsp_src_channel;                                                                            // limiter:rsp_src_channel -> Tiger_MIPS_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                              // Tiger_MIPS_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          addr_router_001_src_endofpacket;                                                                    // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire          addr_router_001_src_valid;                                                                          // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire          addr_router_001_src_startofpacket;                                                                  // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [107:0] addr_router_001_src_data;                                                                           // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire    [4:0] addr_router_001_src_channel;                                                                        // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire          addr_router_001_src_ready;                                                                          // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire          limiter_001_rsp_src_endofpacket;                                                                    // limiter_001:rsp_src_endofpacket -> JTAG_to_FPGA_Bridge_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_001_rsp_src_valid;                                                                          // limiter_001:rsp_src_valid -> JTAG_to_FPGA_Bridge_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_001_rsp_src_startofpacket;                                                                  // limiter_001:rsp_src_startofpacket -> JTAG_to_FPGA_Bridge_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [107:0] limiter_001_rsp_src_data;                                                                           // limiter_001:rsp_src_data -> JTAG_to_FPGA_Bridge_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [4:0] limiter_001_rsp_src_channel;                                                                        // limiter_001:rsp_src_channel -> JTAG_to_FPGA_Bridge_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_001_rsp_src_ready;                                                                          // JTAG_to_FPGA_Bridge_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire          burst_adapter_source0_endofpacket;                                                                  // burst_adapter:source0_endofpacket -> SDRAM_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                        // burst_adapter:source0_valid -> SDRAM_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                // burst_adapter:source0_startofpacket -> SDRAM_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [89:0] burst_adapter_source0_data;                                                                         // burst_adapter:source0_data -> SDRAM_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                        // SDRAM_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire    [4:0] burst_adapter_source0_channel;                                                                      // burst_adapter:source0_channel -> SDRAM_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                     // rst_controller:reset_out -> [Tiger_MIPS:reset, Tiger_MIPS_data_master_translator:reset, Tiger_MIPS_data_master_translator_avalon_universal_master_0_agent:reset, addr_router:reset, cmd_xbar_demux:reset, limiter:reset, rsp_xbar_mux:reset]
	wire          leap_profiler_leap_processor_reset_reset;                                                           // Leap_Profiler:tiger_soft_reset -> rst_controller:reset_in1
	wire          rst_controller_001_reset_out_reset;                                                                 // rst_controller_001:reset_out -> [DCache:reset, DCache_cache_master_translator:reset, DCache_cache_master_translator_avalon_universal_master_0_agent:reset, DCache_cache_slave_translator:reset, DCache_cache_slave_translator_avalon_universal_slave_0_agent:reset, DCache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, JTAG_UART:rst_n, JTAG_UART_avalon_jtag_slave_translator:reset, JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, JTAG_to_FPGA_Bridge_master_translator:reset, JTAG_to_FPGA_Bridge_master_translator_avalon_universal_master_0_agent:reset, Leap_Profiler:reset, Leap_Profiler_leapslave_translator:reset, Leap_Profiler_to_memory_translator:reset, Leap_Sim_Control:reset, Leap_Sim_Control_bridge_master_translator:reset, Leap_Sim_Control_bridge_slave_translator:reset, Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:reset, Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SDRAM:reset_n, SDRAM_s1_translator:reset, SDRAM_s1_translator_avalon_universal_slave_0_agent:reset, SDRAM_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, SDRAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, Tiger_ICache:reset_n, Tiger_ICache_icache_master_translator:reset, Tiger_ICache_icache_master_translator_avalon_universal_master_0_agent:reset, Tiger_ICache_icache_slave_translator:reset, UART:reset_n, UART_s1_translator:reset, UART_s1_translator_avalon_universal_slave_0_agent:reset, UART_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, burst_adapter:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_004:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, limiter_001:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_mux_001:reset, width_adapter:reset, width_adapter_001:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                    // cmd_xbar_demux:src0_endofpacket -> DCache_cache_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                          // cmd_xbar_demux:src0_valid -> DCache_cache_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                  // cmd_xbar_demux:src0_startofpacket -> DCache_cache_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [107:0] cmd_xbar_demux_src0_data;                                                                           // cmd_xbar_demux:src0_data -> DCache_cache_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [4:0] cmd_xbar_demux_src0_channel;                                                                        // cmd_xbar_demux:src0_channel -> DCache_cache_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_src1_endofpacket;                                                                    // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                          // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                  // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [107:0] cmd_xbar_demux_src1_data;                                                                           // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire    [4:0] cmd_xbar_demux_src1_channel;                                                                        // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                          // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_src2_endofpacket;                                                                    // cmd_xbar_demux:src2_endofpacket -> UART_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                          // cmd_xbar_demux:src2_valid -> UART_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                  // cmd_xbar_demux:src2_startofpacket -> UART_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [107:0] cmd_xbar_demux_src2_data;                                                                           // cmd_xbar_demux:src2_data -> UART_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [4:0] cmd_xbar_demux_src2_channel;                                                                        // cmd_xbar_demux:src2_channel -> UART_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                      // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                              // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [107:0] cmd_xbar_demux_001_src0_data;                                                                       // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux_001:sink1_data
	wire    [4:0] cmd_xbar_demux_001_src0_channel;                                                                    // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                      // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                // cmd_xbar_demux_001:src1_endofpacket -> Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                      // cmd_xbar_demux_001:src1_valid -> Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                              // cmd_xbar_demux_001:src1_startofpacket -> Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [107:0] cmd_xbar_demux_001_src1_data;                                                                       // cmd_xbar_demux_001:src1_data -> Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [4:0] cmd_xbar_demux_001_src1_channel;                                                                    // cmd_xbar_demux_001:src1_channel -> Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                      // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_004:sink0_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                              // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	wire  [107:0] cmd_xbar_demux_001_src2_data;                                                                       // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_004:sink0_data
	wire    [4:0] cmd_xbar_demux_001_src2_channel;                                                                    // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_004:sink0_channel
	wire          cmd_xbar_demux_001_src2_ready;                                                                      // cmd_xbar_mux_004:sink0_ready -> cmd_xbar_demux_001:src2_ready
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                                // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                      // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_004:sink1_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                              // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	wire  [107:0] cmd_xbar_demux_002_src0_data;                                                                       // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_004:sink1_data
	wire    [4:0] cmd_xbar_demux_002_src0_channel;                                                                    // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_004:sink1_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                      // cmd_xbar_mux_004:sink1_ready -> cmd_xbar_demux_002:src0_ready
	wire          cmd_xbar_demux_003_src0_endofpacket;                                                                // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_004:sink2_endofpacket
	wire          cmd_xbar_demux_003_src0_valid;                                                                      // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_004:sink2_valid
	wire          cmd_xbar_demux_003_src0_startofpacket;                                                              // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_004:sink2_startofpacket
	wire  [107:0] cmd_xbar_demux_003_src0_data;                                                                       // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_004:sink2_data
	wire    [4:0] cmd_xbar_demux_003_src0_channel;                                                                    // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_004:sink2_channel
	wire          cmd_xbar_demux_003_src0_ready;                                                                      // cmd_xbar_mux_004:sink2_ready -> cmd_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_src0_endofpacket;                                                                    // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                          // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                  // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [107:0] rsp_xbar_demux_src0_data;                                                                           // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire    [4:0] rsp_xbar_demux_src0_channel;                                                                        // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                          // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                      // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                              // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [107:0] rsp_xbar_demux_001_src0_data;                                                                       // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire    [4:0] rsp_xbar_demux_001_src0_channel;                                                                    // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                      // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                                // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                      // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                              // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [107:0] rsp_xbar_demux_001_src1_data;                                                                       // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink0_data
	wire    [4:0] rsp_xbar_demux_001_src1_channel;                                                                    // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                      // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                      // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                              // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [107:0] rsp_xbar_demux_002_src0_data;                                                                       // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire    [4:0] rsp_xbar_demux_002_src0_channel;                                                                    // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                      // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                      // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                              // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [107:0] rsp_xbar_demux_003_src0_data;                                                                       // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink1_data
	wire    [4:0] rsp_xbar_demux_003_src0_channel;                                                                    // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                      // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                      // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                              // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [107:0] rsp_xbar_demux_004_src0_data;                                                                       // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink2_data
	wire    [4:0] rsp_xbar_demux_004_src0_channel;                                                                    // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                      // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_004_src1_endofpacket;                                                                // rsp_xbar_demux_004:src1_endofpacket -> Tiger_ICache_icache_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_004_src1_valid;                                                                      // rsp_xbar_demux_004:src1_valid -> Tiger_ICache_icache_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_004_src1_startofpacket;                                                              // rsp_xbar_demux_004:src1_startofpacket -> Tiger_ICache_icache_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [107:0] rsp_xbar_demux_004_src1_data;                                                                       // rsp_xbar_demux_004:src1_data -> Tiger_ICache_icache_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [4:0] rsp_xbar_demux_004_src1_channel;                                                                    // rsp_xbar_demux_004:src1_channel -> Tiger_ICache_icache_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_004_src2_endofpacket;                                                                // rsp_xbar_demux_004:src2_endofpacket -> DCache_cache_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_004_src2_valid;                                                                      // rsp_xbar_demux_004:src2_valid -> DCache_cache_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_004_src2_startofpacket;                                                              // rsp_xbar_demux_004:src2_startofpacket -> DCache_cache_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [107:0] rsp_xbar_demux_004_src2_data;                                                                       // rsp_xbar_demux_004:src2_data -> DCache_cache_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [4:0] rsp_xbar_demux_004_src2_channel;                                                                    // rsp_xbar_demux_004:src2_channel -> DCache_cache_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_cmd_src_endofpacket;                                                                        // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                      // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [107:0] limiter_cmd_src_data;                                                                               // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire    [4:0] limiter_cmd_src_channel;                                                                            // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_cmd_src_ready;                                                                              // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                       // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                             // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                     // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [107:0] rsp_xbar_mux_src_data;                                                                              // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire    [4:0] rsp_xbar_mux_src_channel;                                                                           // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_src_ready;                                                                             // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire          limiter_001_cmd_src_endofpacket;                                                                    // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          limiter_001_cmd_src_startofpacket;                                                                  // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [107:0] limiter_001_cmd_src_data;                                                                           // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire    [4:0] limiter_001_cmd_src_channel;                                                                        // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire          limiter_001_cmd_src_ready;                                                                          // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                   // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                         // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                 // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [107:0] rsp_xbar_mux_001_src_data;                                                                          // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire    [4:0] rsp_xbar_mux_001_src_channel;                                                                       // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                         // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire          addr_router_002_src_endofpacket;                                                                    // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          addr_router_002_src_valid;                                                                          // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire          addr_router_002_src_startofpacket;                                                                  // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [107:0] addr_router_002_src_data;                                                                           // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire    [4:0] addr_router_002_src_channel;                                                                        // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire          addr_router_002_src_ready;                                                                          // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire          rsp_xbar_demux_004_src1_ready;                                                                      // Tiger_ICache_icache_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_004:src1_ready
	wire          addr_router_003_src_endofpacket;                                                                    // addr_router_003:src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire          addr_router_003_src_valid;                                                                          // addr_router_003:src_valid -> cmd_xbar_demux_003:sink_valid
	wire          addr_router_003_src_startofpacket;                                                                  // addr_router_003:src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire  [107:0] addr_router_003_src_data;                                                                           // addr_router_003:src_data -> cmd_xbar_demux_003:sink_data
	wire    [4:0] addr_router_003_src_channel;                                                                        // addr_router_003:src_channel -> cmd_xbar_demux_003:sink_channel
	wire          addr_router_003_src_ready;                                                                          // cmd_xbar_demux_003:sink_ready -> addr_router_003:src_ready
	wire          rsp_xbar_demux_004_src2_ready;                                                                      // DCache_cache_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_004:src2_ready
	wire          cmd_xbar_demux_src0_ready;                                                                          // DCache_cache_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src0_ready
	wire          id_router_src_endofpacket;                                                                          // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                        // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [107:0] id_router_src_data;                                                                                 // id_router:src_data -> rsp_xbar_demux:sink_data
	wire    [4:0] id_router_src_channel;                                                                              // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                   // cmd_xbar_mux_001:src_endofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                         // cmd_xbar_mux_001:src_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                 // cmd_xbar_mux_001:src_startofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [107:0] cmd_xbar_mux_001_src_data;                                                                          // cmd_xbar_mux_001:src_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [4:0] cmd_xbar_mux_001_src_channel;                                                                       // cmd_xbar_mux_001:src_channel -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                         // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire          id_router_001_src_endofpacket;                                                                      // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                            // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                    // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [107:0] id_router_001_src_data;                                                                             // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire    [4:0] id_router_001_src_channel;                                                                          // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                            // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_demux_src2_ready;                                                                          // UART_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src2_ready
	wire          id_router_002_src_endofpacket;                                                                      // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                            // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                    // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [107:0] id_router_002_src_data;                                                                             // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire    [4:0] id_router_002_src_channel;                                                                          // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                            // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_demux_001_src1_ready;                                                                      // Leap_Sim_Control_bridge_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src1_ready
	wire          id_router_003_src_endofpacket;                                                                      // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                            // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                    // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [107:0] id_router_003_src_data;                                                                             // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire    [4:0] id_router_003_src_channel;                                                                          // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                            // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_mux_004_src_endofpacket;                                                                   // cmd_xbar_mux_004:src_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_mux_004_src_valid;                                                                         // cmd_xbar_mux_004:src_valid -> width_adapter:in_valid
	wire          cmd_xbar_mux_004_src_startofpacket;                                                                 // cmd_xbar_mux_004:src_startofpacket -> width_adapter:in_startofpacket
	wire  [107:0] cmd_xbar_mux_004_src_data;                                                                          // cmd_xbar_mux_004:src_data -> width_adapter:in_data
	wire    [4:0] cmd_xbar_mux_004_src_channel;                                                                       // cmd_xbar_mux_004:src_channel -> width_adapter:in_channel
	wire          cmd_xbar_mux_004_src_ready;                                                                         // width_adapter:in_ready -> cmd_xbar_mux_004:src_ready
	wire          width_adapter_src_endofpacket;                                                                      // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                            // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                    // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [89:0] width_adapter_src_data;                                                                             // width_adapter:out_data -> burst_adapter:sink0_data
	wire          width_adapter_src_ready;                                                                            // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire    [4:0] width_adapter_src_channel;                                                                          // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire          id_router_004_src_endofpacket;                                                                      // id_router_004:src_endofpacket -> width_adapter_001:in_endofpacket
	wire          id_router_004_src_valid;                                                                            // id_router_004:src_valid -> width_adapter_001:in_valid
	wire          id_router_004_src_startofpacket;                                                                    // id_router_004:src_startofpacket -> width_adapter_001:in_startofpacket
	wire   [89:0] id_router_004_src_data;                                                                             // id_router_004:src_data -> width_adapter_001:in_data
	wire    [4:0] id_router_004_src_channel;                                                                          // id_router_004:src_channel -> width_adapter_001:in_channel
	wire          id_router_004_src_ready;                                                                            // width_adapter_001:in_ready -> id_router_004:src_ready
	wire          width_adapter_001_src_endofpacket;                                                                  // width_adapter_001:out_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          width_adapter_001_src_valid;                                                                        // width_adapter_001:out_valid -> rsp_xbar_demux_004:sink_valid
	wire          width_adapter_001_src_startofpacket;                                                                // width_adapter_001:out_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [107:0] width_adapter_001_src_data;                                                                         // width_adapter_001:out_data -> rsp_xbar_demux_004:sink_data
	wire          width_adapter_001_src_ready;                                                                        // rsp_xbar_demux_004:sink_ready -> width_adapter_001:out_ready
	wire    [4:0] width_adapter_001_src_channel;                                                                      // width_adapter_001:out_channel -> rsp_xbar_demux_004:sink_channel
	wire    [4:0] limiter_cmd_valid_data;                                                                             // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire    [4:0] limiter_001_cmd_valid_data;                                                                         // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid

	tiger_top #(
		.RESET_ADDRESS (1073741824)
	) tiger_mips (
		.clk                           (clk_clk),                                     //              clock.clk
		.reset                         (rst_controller_reset_out_reset),              //              reset.reset
		.avm_instrMaster_address       (tiger_mips_instruction_master_address),       // instruction_master.address
		.avm_instrMaster_read          (tiger_mips_instruction_master_read),          //                   .read
		.avm_instrMaster_write         (tiger_mips_instruction_master_write),         //                   .write
		.avm_instrMaster_writedata     (tiger_mips_instruction_master_writedata),     //                   .writedata
		.avm_instrMaster_byteenable    (tiger_mips_instruction_master_byteenable),    //                   .byteenable
		.avm_instrMaster_readdata      (tiger_mips_instruction_master_readdata),      //                   .readdata
		.avm_instrMaster_waitrequest   (tiger_mips_instruction_master_waitrequest),   //                   .waitrequest
		.avm_instrMaster_readdatavalid (tiger_mips_instruction_master_readdatavalid), //                   .readdatavalid
		.avm_dataMaster_address        (tiger_mips_data_master_address),              //        data_master.address
		.avm_dataMaster_read           (tiger_mips_data_master_read),                 //                   .read
		.avm_dataMaster_write          (tiger_mips_data_master_write),                //                   .write
		.avm_dataMaster_writedata      (tiger_mips_data_master_writedata),            //                   .writedata
		.avm_dataMaster_byteenable     (tiger_mips_data_master_byteenable),           //                   .byteenable
		.avm_dataMaster_readdata       (tiger_mips_data_master_readdata),             //                   .readdata
		.avm_dataMaster_waitrequest    (tiger_mips_data_master_waitrequest),          //                   .waitrequest
		.avm_dataMaster_readdatavalid  (tiger_mips_data_master_readdatavalid)         //                   .readdatavalid
	);

	LeapTop #(
		.STARTING_PC   (1073741856),
		.prof_param_N2 (8),
		.prof_param_S2 (5),
		.prof_param_CW (32)
	) leap_profiler (
		.clk                         (clk_clk),                                                          //                clock.clk
		.reset                       (rst_controller_001_reset_out_reset),                               //                reset.reset
		.tiger_soft_reset            (leap_profiler_leap_processor_reset_reset),                         // leap_processor_reset.reset
		.avs_from_cpu_address        (tiger_mips_instruction_master_address),                            //             from_cpu.address
		.avs_from_cpu_read           (tiger_mips_instruction_master_read),                               //                     .read
		.avs_from_cpu_write          (tiger_mips_instruction_master_write),                              //                     .write
		.avs_from_cpu_writedata      (tiger_mips_instruction_master_writedata),                          //                     .writedata
		.avs_from_cpu_byteenable     (tiger_mips_instruction_master_byteenable),                         //                     .byteenable
		.avs_from_cpu_readdata       (tiger_mips_instruction_master_readdata),                           //                     .readdata
		.avs_from_cpu_waitrequest    (tiger_mips_instruction_master_waitrequest),                        //                     .waitrequest
		.avs_from_cpu_readdatavalid  (tiger_mips_instruction_master_readdatavalid),                      //                     .readdatavalid
		.avs_to_memory_address       (leap_profiler_to_memory_address),                                  //            to_memory.address
		.avs_to_memory_read          (leap_profiler_to_memory_read),                                     //                     .read
		.avs_to_memory_write         (leap_profiler_to_memory_write),                                    //                     .write
		.avs_to_memory_writedata     (leap_profiler_to_memory_writedata),                                //                     .writedata
		.avs_to_memory_byteenable    (leap_profiler_to_memory_byteenable),                               //                     .byteenable
		.avs_to_memory_readdata      (leap_profiler_to_memory_readdata),                                 //                     .readdata
		.avs_to_memory_waitrequest   (leap_profiler_to_memory_waitrequest),                              //                     .waitrequest
		.avs_to_memory_readdatavalid (leap_profiler_to_memory_readdatavalid),                            //                     .readdatavalid
		.avs_leapSlave_address       (leap_profiler_leapslave_translator_avalon_anti_slave_0_address),   //            leapslave.address
		.avs_leapSlave_read          (leap_profiler_leapslave_translator_avalon_anti_slave_0_read),      //                     .read
		.avs_leapSlave_write         (leap_profiler_leapslave_translator_avalon_anti_slave_0_write),     //                     .write
		.avs_leapSlave_writedata     (leap_profiler_leapslave_translator_avalon_anti_slave_0_writedata), //                     .writedata
		.avs_leapSlave_readdata      (leap_profiler_leapslave_translator_avalon_anti_slave_0_readdata),  //                     .readdata
		.coe_exe_start               (leap_profiling_signals_start),                                     //    profiling_signals.export
		.coe_exe_end                 (leap_profiling_signals_end),                                       //                     .export
		.coe_debug_select            (leap_debug_port_select),                                           //           debug_port.export
		.coe_debug_lights            (leap_debug_port_lights)                                            //                     .export
	);

	leap_sim_controller #(
		.STARTING_PC (1073741856),
		.N2          (8)
	) leap_sim_control (
		.clk                           (clk_clk),                                                                //         clock.clk
		.reset                         (rst_controller_001_reset_out_reset),                                     //         reset.reset
		.avs_bridge_slave_address      (leap_sim_control_bridge_slave_translator_avalon_anti_slave_0_address),   //  bridge_slave.address
		.avs_bridge_slave_read         (leap_sim_control_bridge_slave_translator_avalon_anti_slave_0_read),      //              .read
		.avs_bridge_slave_write        (leap_sim_control_bridge_slave_translator_avalon_anti_slave_0_write),     //              .write
		.avs_bridge_slave_writedata    (leap_sim_control_bridge_slave_translator_avalon_anti_slave_0_writedata), //              .writedata
		.avs_bridge_slave_readdata     (leap_sim_control_bridge_slave_translator_avalon_anti_slave_0_readdata),  //              .readdata
		.avm_bridge_master_readdata    (leap_sim_control_bridge_master_readdata),                                // bridge_master.readdata
		.avm_bridge_master_waitrequest (leap_sim_control_bridge_master_waitrequest),                             //              .waitrequest
		.avm_bridge_master_address     (leap_sim_control_bridge_master_address),                                 //              .address
		.avm_bridge_master_byteenable  (leap_sim_control_bridge_master_byteenable),                              //              .byteenable
		.avm_bridge_master_read        (leap_sim_control_bridge_master_read),                                    //              .read
		.avm_bridge_master_write       (leap_sim_control_bridge_master_write),                                   //              .write
		.avm_bridge_master_writedata   (leap_sim_control_bridge_master_writedata)                                //              .writedata
	);

	tiger_icache_av_1port tiger_icache (
		.clk                                  (clk_clk),                                                                //         clock.clk
		.reset_n                              (~rst_controller_001_reset_out_reset),                                    //         reset.reset_n
		.avs_icache_slave_address             (tiger_icache_icache_slave_translator_avalon_anti_slave_0_address),       //  icache_slave.address
		.avs_icache_slave_read                (tiger_icache_icache_slave_translator_avalon_anti_slave_0_read),          //              .read
		.avs_icache_slave_readdata            (tiger_icache_icache_slave_translator_avalon_anti_slave_0_readdata),      //              .readdata
		.avs_icache_slave_readdatavalid       (tiger_icache_icache_slave_translator_avalon_anti_slave_0_readdatavalid), //              .readdatavalid
		.avs_icache_slave_waitrequest         (tiger_icache_icache_slave_translator_avalon_anti_slave_0_waitrequest),   //              .waitrequest
		.avm_icache_master_readdata           (tiger_icache_icache_master_readdata),                                    // icache_master.readdata
		.avm_icache_master_readdatavalid      (tiger_icache_icache_master_readdatavalid),                               //              .readdatavalid
		.avm_icache_master_waitrequest        (tiger_icache_icache_master_waitrequest),                                 //              .waitrequest
		.avm_icache_master_address            (tiger_icache_icache_master_address),                                     //              .address
		.avm_icache_master_beginbursttransfer (tiger_icache_icache_master_beginbursttransfer),                          //              .beginbursttransfer
		.avm_icache_master_burstcount         (tiger_icache_icache_master_burstcount),                                  //              .burstcount
		.avm_icache_master_read               (tiger_icache_icache_master_read)                                         //              .read
	);

	legup_dm_wt_cache dcache (
		.reset                   (rst_controller_001_reset_out_reset),                              //        reset.reset
		.clk                     (clk_clk),                                                         //          clk.clk
		.avs_cache_address       (dcache_cache_slave_translator_avalon_anti_slave_0_address),       //  cache_slave.address
		.avs_cache_byteenable    (dcache_cache_slave_translator_avalon_anti_slave_0_byteenable),    //             .byteenable
		.avs_cache_read          (dcache_cache_slave_translator_avalon_anti_slave_0_read),          //             .read
		.avs_cache_write         (dcache_cache_slave_translator_avalon_anti_slave_0_write),         //             .write
		.avs_cache_writedata     (dcache_cache_slave_translator_avalon_anti_slave_0_writedata),     //             .writedata
		.avs_cache_readdata      (dcache_cache_slave_translator_avalon_anti_slave_0_readdata),      //             .readdata
		.avs_cache_readdatavalid (dcache_cache_slave_translator_avalon_anti_slave_0_readdatavalid), //             .readdatavalid
		.avs_cache_waitrequest   (dcache_cache_slave_translator_avalon_anti_slave_0_waitrequest),   //             .waitrequest
		.avm_cache_readdata      (dcache_cache_master_readdata),                                    // cache_master.readdata
		.avm_cache_readdatavalid (dcache_cache_master_readdatavalid),                               //             .readdatavalid
		.avm_cache_waitrequest   (dcache_cache_master_waitrequest),                                 //             .waitrequest
		.avm_cache_address       (dcache_cache_master_address),                                     //             .address
		.avm_cache_burstcount    (dcache_cache_master_burstcount),                                  //             .burstcount
		.avm_cache_byteenable    (dcache_cache_master_byteenable),                                  //             .byteenable
		.avm_cache_read          (dcache_cache_master_read),                                        //             .read
		.avm_cache_write         (dcache_cache_master_write),                                       //             .write
		.avm_cache_writedata     (dcache_cache_master_writedata)                                    //             .writedata
	);

	legup_system_JTAG_to_FPGA_Bridge #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) jtag_to_fpga_bridge (
		.clk_clk              (clk_clk),                                  //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                           //    clk_reset.reset
		.master_address       (jtag_to_fpga_bridge_master_address),       //       master.address
		.master_readdata      (jtag_to_fpga_bridge_master_readdata),      //             .readdata
		.master_read          (jtag_to_fpga_bridge_master_read),          //             .read
		.master_write         (jtag_to_fpga_bridge_master_write),         //             .write
		.master_writedata     (jtag_to_fpga_bridge_master_writedata),     //             .writedata
		.master_waitrequest   (jtag_to_fpga_bridge_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (jtag_to_fpga_bridge_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (jtag_to_fpga_bridge_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                          // master_reset.reset
	);

	legup_system_SDRAM sdram (
		.clk            (clk_clk),                                               //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                   // reset.reset_n
		.az_addr        (sdram_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                                       //  wire.export
		.zs_ba          (sdram_wire_ba),                                         //      .export
		.zs_cas_n       (sdram_wire_cas_n),                                      //      .export
		.zs_cke         (sdram_wire_cke),                                        //      .export
		.zs_cs_n        (sdram_wire_cs_n),                                       //      .export
		.zs_dq          (sdram_wire_dq),                                         //      .export
		.zs_dqm         (sdram_wire_dqm),                                        //      .export
		.zs_ras_n       (sdram_wire_ras_n),                                      //      .export
		.zs_we_n        (sdram_wire_we_n)                                        //      .export
	);

	legup_system_JTAG_UART jtag_uart (
		.clk            (clk_clk),                                                                //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                                    //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         ()                                                                        //               irq.irq
	);

	legup_system_UART uart (
		.clk           (clk_clk),                                              //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                  //               reset.reset_n
		.address       (uart_s1_translator_avalon_anti_slave_0_address),       //                  s1.address
		.begintransfer (uart_s1_translator_avalon_anti_slave_0_begintransfer), //                    .begintransfer
		.chipselect    (uart_s1_translator_avalon_anti_slave_0_chipselect),    //                    .chipselect
		.read_n        (~uart_s1_translator_avalon_anti_slave_0_read),         //                    .read_n
		.write_n       (~uart_s1_translator_avalon_anti_slave_0_write),        //                    .write_n
		.writedata     (uart_s1_translator_avalon_anti_slave_0_writedata),     //                    .writedata
		.readdata      (uart_s1_translator_avalon_anti_slave_0_readdata),      //                    .readdata
		.dataavailable (),                                                     //                    .dataavailable
		.readyfordata  (),                                                     //                    .readyfordata
		.rxd           (uart_wire_rxd),                                        // external_connection.export
		.txd           (uart_wire_txd),                                        //                    .export
		.irq           ()                                                      //                 irq.irq
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) leap_sim_control_bridge_master_translator (
		.clk                      (clk_clk),                                                                           //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                //                     reset.reset
		.uav_address              (leap_sim_control_bridge_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (leap_sim_control_bridge_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (leap_sim_control_bridge_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (leap_sim_control_bridge_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (leap_sim_control_bridge_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (leap_sim_control_bridge_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (leap_sim_control_bridge_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (leap_sim_control_bridge_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (leap_sim_control_bridge_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (leap_sim_control_bridge_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (leap_sim_control_bridge_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (leap_sim_control_bridge_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (leap_sim_control_bridge_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (leap_sim_control_bridge_master_byteenable),                                         //                          .byteenable
		.av_read                  (leap_sim_control_bridge_master_read),                                               //                          .read
		.av_readdata              (leap_sim_control_bridge_master_readdata),                                           //                          .readdata
		.av_write                 (leap_sim_control_bridge_master_write),                                              //                          .write
		.av_writedata             (leap_sim_control_bridge_master_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                              //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                              //               (terminated)
		.av_begintransfer         (1'b0),                                                                              //               (terminated)
		.av_chipselect            (1'b0),                                                                              //               (terminated)
		.av_readdatavalid         (),                                                                                  //               (terminated)
		.av_lock                  (1'b0),                                                                              //               (terminated)
		.av_debugaccess           (1'b0),                                                                              //               (terminated)
		.uav_clken                (),                                                                                  //               (terminated)
		.av_clken                 (1'b1),                                                                              //               (terminated)
		.uav_response             (2'b00),                                                                             //               (terminated)
		.av_response              (),                                                                                  //               (terminated)
		.uav_writeresponserequest (),                                                                                  //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                              //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                              //               (terminated)
		.av_writeresponsevalid    ()                                                                                   //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (30),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) leap_profiler_leapslave_translator (
		.clk                      (clk_clk),                                                                           //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                //                    reset.reset
		.uav_address              (leap_sim_control_bridge_master_translator_avalon_universal_master_0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (leap_sim_control_bridge_master_translator_avalon_universal_master_0_burstcount),    //                         .burstcount
		.uav_read                 (leap_sim_control_bridge_master_translator_avalon_universal_master_0_read),          //                         .read
		.uav_write                (leap_sim_control_bridge_master_translator_avalon_universal_master_0_write),         //                         .write
		.uav_waitrequest          (leap_sim_control_bridge_master_translator_avalon_universal_master_0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (leap_sim_control_bridge_master_translator_avalon_universal_master_0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (leap_sim_control_bridge_master_translator_avalon_universal_master_0_byteenable),    //                         .byteenable
		.uav_readdata             (leap_sim_control_bridge_master_translator_avalon_universal_master_0_readdata),      //                         .readdata
		.uav_writedata            (leap_sim_control_bridge_master_translator_avalon_universal_master_0_writedata),     //                         .writedata
		.uav_lock                 (leap_sim_control_bridge_master_translator_avalon_universal_master_0_lock),          //                         .lock
		.uav_debugaccess          (leap_sim_control_bridge_master_translator_avalon_universal_master_0_debugaccess),   //                         .debugaccess
		.av_address               (leap_profiler_leapslave_translator_avalon_anti_slave_0_address),                    //      avalon_anti_slave_0.address
		.av_write                 (leap_profiler_leapslave_translator_avalon_anti_slave_0_write),                      //                         .write
		.av_read                  (leap_profiler_leapslave_translator_avalon_anti_slave_0_read),                       //                         .read
		.av_readdata              (leap_profiler_leapslave_translator_avalon_anti_slave_0_readdata),                   //                         .readdata
		.av_writedata             (leap_profiler_leapslave_translator_avalon_anti_slave_0_writedata),                  //                         .writedata
		.av_begintransfer         (),                                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                                  //              (terminated)
		.av_burstcount            (),                                                                                  //              (terminated)
		.av_byteenable            (),                                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                                              //              (terminated)
		.av_writebyteenable       (),                                                                                  //              (terminated)
		.av_lock                  (),                                                                                  //              (terminated)
		.av_chipselect            (),                                                                                  //              (terminated)
		.av_clken                 (),                                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                                              //              (terminated)
		.av_debugaccess           (),                                                                                  //              (terminated)
		.av_outputenable          (),                                                                                  //              (terminated)
		.uav_response             (),                                                                                  //              (terminated)
		.av_response              (2'b00),                                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                               //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) leap_profiler_to_memory_translator (
		.clk                      (clk_clk),                                                                    //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                         //                     reset.reset
		.uav_address              (leap_profiler_to_memory_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (leap_profiler_to_memory_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (leap_profiler_to_memory_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (leap_profiler_to_memory_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (leap_profiler_to_memory_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (leap_profiler_to_memory_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (leap_profiler_to_memory_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (leap_profiler_to_memory_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (leap_profiler_to_memory_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (leap_profiler_to_memory_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (leap_profiler_to_memory_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (leap_profiler_to_memory_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (leap_profiler_to_memory_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (leap_profiler_to_memory_byteenable),                                         //                          .byteenable
		.av_read                  (leap_profiler_to_memory_read),                                               //                          .read
		.av_readdata              (leap_profiler_to_memory_readdata),                                           //                          .readdata
		.av_readdatavalid         (leap_profiler_to_memory_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (leap_profiler_to_memory_write),                                              //                          .write
		.av_writedata             (leap_profiler_to_memory_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                       //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                       //               (terminated)
		.av_begintransfer         (1'b0),                                                                       //               (terminated)
		.av_chipselect            (1'b0),                                                                       //               (terminated)
		.av_lock                  (1'b0),                                                                       //               (terminated)
		.av_debugaccess           (1'b0),                                                                       //               (terminated)
		.uav_clken                (),                                                                           //               (terminated)
		.av_clken                 (1'b1),                                                                       //               (terminated)
		.uav_response             (2'b00),                                                                      //               (terminated)
		.av_response              (),                                                                           //               (terminated)
		.uav_writeresponserequest (),                                                                           //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                       //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                       //               (terminated)
		.av_writeresponsevalid    ()                                                                            //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (30),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) tiger_icache_icache_slave_translator (
		.clk                      (clk_clk),                                                                    //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                         //                    reset.reset
		.uav_address              (leap_profiler_to_memory_translator_avalon_universal_master_0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (leap_profiler_to_memory_translator_avalon_universal_master_0_burstcount),    //                         .burstcount
		.uav_read                 (leap_profiler_to_memory_translator_avalon_universal_master_0_read),          //                         .read
		.uav_write                (leap_profiler_to_memory_translator_avalon_universal_master_0_write),         //                         .write
		.uav_waitrequest          (leap_profiler_to_memory_translator_avalon_universal_master_0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (leap_profiler_to_memory_translator_avalon_universal_master_0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (leap_profiler_to_memory_translator_avalon_universal_master_0_byteenable),    //                         .byteenable
		.uav_readdata             (leap_profiler_to_memory_translator_avalon_universal_master_0_readdata),      //                         .readdata
		.uav_writedata            (leap_profiler_to_memory_translator_avalon_universal_master_0_writedata),     //                         .writedata
		.uav_lock                 (leap_profiler_to_memory_translator_avalon_universal_master_0_lock),          //                         .lock
		.uav_debugaccess          (leap_profiler_to_memory_translator_avalon_universal_master_0_debugaccess),   //                         .debugaccess
		.av_address               (tiger_icache_icache_slave_translator_avalon_anti_slave_0_address),           //      avalon_anti_slave_0.address
		.av_read                  (tiger_icache_icache_slave_translator_avalon_anti_slave_0_read),              //                         .read
		.av_readdata              (tiger_icache_icache_slave_translator_avalon_anti_slave_0_readdata),          //                         .readdata
		.av_readdatavalid         (tiger_icache_icache_slave_translator_avalon_anti_slave_0_readdatavalid),     //                         .readdatavalid
		.av_waitrequest           (tiger_icache_icache_slave_translator_avalon_anti_slave_0_waitrequest),       //                         .waitrequest
		.av_write                 (),                                                                           //              (terminated)
		.av_writedata             (),                                                                           //              (terminated)
		.av_begintransfer         (),                                                                           //              (terminated)
		.av_beginbursttransfer    (),                                                                           //              (terminated)
		.av_burstcount            (),                                                                           //              (terminated)
		.av_byteenable            (),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                           //              (terminated)
		.av_lock                  (),                                                                           //              (terminated)
		.av_chipselect            (),                                                                           //              (terminated)
		.av_clken                 (),                                                                           //              (terminated)
		.uav_clken                (1'b0),                                                                       //              (terminated)
		.av_debugaccess           (),                                                                           //              (terminated)
		.av_outputenable          (),                                                                           //              (terminated)
		.uav_response             (),                                                                           //              (terminated)
		.av_response              (2'b00),                                                                      //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                       //              (terminated)
		.uav_writeresponsevalid   (),                                                                           //              (terminated)
		.av_writeresponserequest  (),                                                                           //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                        //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) tiger_mips_data_master_translator (
		.clk                      (clk_clk),                                                                   //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                            //                     reset.reset
		.uav_address              (tiger_mips_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (tiger_mips_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (tiger_mips_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (tiger_mips_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (tiger_mips_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (tiger_mips_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (tiger_mips_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (tiger_mips_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (tiger_mips_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (tiger_mips_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (tiger_mips_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (tiger_mips_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (tiger_mips_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (tiger_mips_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (tiger_mips_data_master_read),                                               //                          .read
		.av_readdata              (tiger_mips_data_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (tiger_mips_data_master_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (tiger_mips_data_master_write),                                              //                          .write
		.av_writedata             (tiger_mips_data_master_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                      //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                      //               (terminated)
		.av_begintransfer         (1'b0),                                                                      //               (terminated)
		.av_chipselect            (1'b0),                                                                      //               (terminated)
		.av_lock                  (1'b0),                                                                      //               (terminated)
		.av_debugaccess           (1'b0),                                                                      //               (terminated)
		.uav_clken                (),                                                                          //               (terminated)
		.av_clken                 (1'b1),                                                                      //               (terminated)
		.uav_response             (2'b00),                                                                     //               (terminated)
		.av_response              (),                                                                          //               (terminated)
		.uav_writeresponserequest (),                                                                          //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                      //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                      //               (terminated)
		.av_writeresponsevalid    ()                                                                           //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) jtag_to_fpga_bridge_master_translator (
		.clk                      (clk_clk),                                                                       //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                            //                     reset.reset
		.uav_address              (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (jtag_to_fpga_bridge_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (jtag_to_fpga_bridge_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (jtag_to_fpga_bridge_master_byteenable),                                         //                          .byteenable
		.av_read                  (jtag_to_fpga_bridge_master_read),                                               //                          .read
		.av_readdata              (jtag_to_fpga_bridge_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (jtag_to_fpga_bridge_master_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (jtag_to_fpga_bridge_master_write),                                              //                          .write
		.av_writedata             (jtag_to_fpga_bridge_master_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                          //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                          //               (terminated)
		.av_begintransfer         (1'b0),                                                                          //               (terminated)
		.av_chipselect            (1'b0),                                                                          //               (terminated)
		.av_lock                  (1'b0),                                                                          //               (terminated)
		.av_debugaccess           (1'b0),                                                                          //               (terminated)
		.uav_clken                (),                                                                              //               (terminated)
		.av_clken                 (1'b1),                                                                          //               (terminated)
		.uav_response             (2'b00),                                                                         //               (terminated)
		.av_response              (),                                                                              //               (terminated)
		.uav_writeresponserequest (),                                                                              //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                          //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                          //               (terminated)
		.av_writeresponsevalid    ()                                                                               //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (6),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (8),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (1),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) tiger_icache_icache_master_translator (
		.clk                      (clk_clk),                                                                       //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                            //                     reset.reset
		.uav_address              (tiger_icache_icache_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (tiger_icache_icache_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (tiger_icache_icache_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (tiger_icache_icache_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (tiger_icache_icache_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (tiger_icache_icache_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (tiger_icache_icache_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (tiger_icache_icache_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (tiger_icache_icache_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (tiger_icache_icache_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (tiger_icache_icache_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (tiger_icache_icache_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (tiger_icache_icache_master_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (tiger_icache_icache_master_burstcount),                                         //                          .burstcount
		.av_beginbursttransfer    (tiger_icache_icache_master_beginbursttransfer),                                 //                          .beginbursttransfer
		.av_read                  (tiger_icache_icache_master_read),                                               //                          .read
		.av_readdata              (tiger_icache_icache_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (tiger_icache_icache_master_readdatavalid),                                      //                          .readdatavalid
		.av_byteenable            (4'b1111),                                                                       //               (terminated)
		.av_begintransfer         (1'b0),                                                                          //               (terminated)
		.av_chipselect            (1'b0),                                                                          //               (terminated)
		.av_write                 (1'b0),                                                                          //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                          //               (terminated)
		.av_lock                  (1'b0),                                                                          //               (terminated)
		.av_debugaccess           (1'b0),                                                                          //               (terminated)
		.uav_clken                (),                                                                              //               (terminated)
		.av_clken                 (1'b1),                                                                          //               (terminated)
		.uav_response             (2'b00),                                                                         //               (terminated)
		.av_response              (),                                                                              //               (terminated)
		.uav_writeresponserequest (),                                                                              //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                          //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                          //               (terminated)
		.av_writeresponsevalid    ()                                                                               //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (3),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (5),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) dcache_cache_master_translator (
		.clk                      (clk_clk),                                                                //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                     //                     reset.reset
		.uav_address              (dcache_cache_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (dcache_cache_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (dcache_cache_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (dcache_cache_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (dcache_cache_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (dcache_cache_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (dcache_cache_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (dcache_cache_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (dcache_cache_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (dcache_cache_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (dcache_cache_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (dcache_cache_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (dcache_cache_master_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (dcache_cache_master_burstcount),                                         //                          .burstcount
		.av_byteenable            (dcache_cache_master_byteenable),                                         //                          .byteenable
		.av_read                  (dcache_cache_master_read),                                               //                          .read
		.av_readdata              (dcache_cache_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (dcache_cache_master_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (dcache_cache_master_write),                                              //                          .write
		.av_writedata             (dcache_cache_master_writedata),                                          //                          .writedata
		.av_beginbursttransfer    (1'b0),                                                                   //               (terminated)
		.av_begintransfer         (1'b0),                                                                   //               (terminated)
		.av_chipselect            (1'b0),                                                                   //               (terminated)
		.av_lock                  (1'b0),                                                                   //               (terminated)
		.av_debugaccess           (1'b0),                                                                   //               (terminated)
		.uav_clken                (),                                                                       //               (terminated)
		.av_clken                 (1'b1),                                                                   //               (terminated)
		.uav_response             (2'b00),                                                                  //               (terminated)
		.av_response              (),                                                                       //               (terminated)
		.uav_writeresponserequest (),                                                                       //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                   //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                   //               (terminated)
		.av_writeresponsevalid    ()                                                                        //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (31),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dcache_cache_slave_translator (
		.clk                      (clk_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                            //                    reset.reset
		.uav_address              (dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (dcache_cache_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (dcache_cache_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (dcache_cache_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (dcache_cache_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (dcache_cache_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (dcache_cache_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (dcache_cache_slave_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (dcache_cache_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer         (),                                                                              //              (terminated)
		.av_beginbursttransfer    (),                                                                              //              (terminated)
		.av_burstcount            (),                                                                              //              (terminated)
		.av_writebyteenable       (),                                                                              //              (terminated)
		.av_lock                  (),                                                                              //              (terminated)
		.av_chipselect            (),                                                                              //              (terminated)
		.av_clken                 (),                                                                              //              (terminated)
		.uav_clken                (1'b0),                                                                          //              (terminated)
		.av_debugaccess           (),                                                                              //              (terminated)
		.av_outputenable          (),                                                                              //              (terminated)
		.uav_response             (),                                                                              //              (terminated)
		.av_response              (2'b00),                                                                         //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                          //              (terminated)
		.uav_writeresponsevalid   (),                                                                              //              (terminated)
		.av_writeresponserequest  (),                                                                              //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                      (clk_clk),                                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                     //                    reset.reset
		.uav_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                                       //              (terminated)
		.av_burstcount            (),                                                                                       //              (terminated)
		.av_byteenable            (),                                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                                       //              (terminated)
		.av_lock                  (),                                                                                       //              (terminated)
		.av_clken                 (),                                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                                   //              (terminated)
		.av_debugaccess           (),                                                                                       //              (terminated)
		.av_outputenable          (),                                                                                       //              (terminated)
		.uav_response             (),                                                                                       //              (terminated)
		.av_response              (2'b00),                                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) uart_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                 //                    reset.reset
		.uav_address              (uart_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (uart_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (uart_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (uart_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (uart_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (uart_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (uart_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (uart_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (uart_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (uart_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (uart_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (uart_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (uart_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (uart_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (uart_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (uart_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (uart_s1_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_chipselect            (uart_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (8),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) leap_sim_control_bridge_slave_translator (
		.clk                      (clk_clk),                                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                       //                    reset.reset
		.uav_address              (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (leap_sim_control_bridge_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (leap_sim_control_bridge_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (leap_sim_control_bridge_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (leap_sim_control_bridge_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (leap_sim_control_bridge_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                                         //              (terminated)
		.av_burstcount            (),                                                                                         //              (terminated)
		.av_byteenable            (),                                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                                         //              (terminated)
		.av_lock                  (),                                                                                         //              (terminated)
		.av_chipselect            (),                                                                                         //              (terminated)
		.av_clken                 (),                                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                                     //              (terminated)
		.av_debugaccess           (),                                                                                         //              (terminated)
		.av_outputenable          (),                                                                                         //              (terminated)
		.uav_response             (),                                                                                         //              (terminated)
		.av_response              (2'b00),                                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_s1_translator (
		.clk                      (clk_clk),                                                             //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                  //                    reset.reset
		.uav_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sdram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sdram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sdram_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sdram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sdram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (sdram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (sdram_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (sdram_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (sdram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_BEGIN_BURST           (90),
		.PKT_BURSTWRAP_H           (82),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BURST_SIZE_H          (85),
		.PKT_BURST_SIZE_L          (83),
		.PKT_BURST_TYPE_H          (87),
		.PKT_BURST_TYPE_L          (86),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (92),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (95),
		.PKT_THREAD_ID_H           (98),
		.PKT_THREAD_ID_L           (98),
		.PKT_CACHE_H               (105),
		.PKT_CACHE_L               (102),
		.PKT_DATA_SIDEBAND_H       (89),
		.PKT_DATA_SIDEBAND_L       (89),
		.PKT_QOS_H                 (91),
		.PKT_QOS_L                 (91),
		.PKT_ADDR_SIDEBAND_H       (88),
		.PKT_ADDR_SIDEBAND_L       (88),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_RESPONSE_STATUS_L     (106),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (5),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (3),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) tiger_mips_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                            //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.av_address              (tiger_mips_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (tiger_mips_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (tiger_mips_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (tiger_mips_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (tiger_mips_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (tiger_mips_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (tiger_mips_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (tiger_mips_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (tiger_mips_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (tiger_mips_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (tiger_mips_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (tiger_mips_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (tiger_mips_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (tiger_mips_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (tiger_mips_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (tiger_mips_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_rsp_src_valid),                                                              //        rp.valid
		.rp_data                 (limiter_rsp_src_data),                                                               //          .data
		.rp_channel              (limiter_rsp_src_channel),                                                            //          .channel
		.rp_startofpacket        (limiter_rsp_src_startofpacket),                                                      //          .startofpacket
		.rp_endofpacket          (limiter_rsp_src_endofpacket),                                                        //          .endofpacket
		.rp_ready                (limiter_rsp_src_ready),                                                              //          .ready
		.av_response             (),                                                                                   // (terminated)
		.av_writeresponserequest (1'b0),                                                                               // (terminated)
		.av_writeresponsevalid   ()                                                                                    // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_BEGIN_BURST           (90),
		.PKT_BURSTWRAP_H           (82),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BURST_SIZE_H          (85),
		.PKT_BURST_SIZE_L          (83),
		.PKT_BURST_TYPE_H          (87),
		.PKT_BURST_TYPE_L          (86),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (92),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (95),
		.PKT_THREAD_ID_H           (98),
		.PKT_THREAD_ID_L           (98),
		.PKT_CACHE_H               (105),
		.PKT_CACHE_L               (102),
		.PKT_DATA_SIDEBAND_H       (89),
		.PKT_DATA_SIDEBAND_L       (89),
		.PKT_QOS_H                 (91),
		.PKT_QOS_L                 (91),
		.PKT_ADDR_SIDEBAND_H       (88),
		.PKT_ADDR_SIDEBAND_L       (88),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_RESPONSE_STATUS_L     (106),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (5),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                                //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.av_address              (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_001_rsp_src_valid),                                                              //        rp.valid
		.rp_data                 (limiter_001_rsp_src_data),                                                               //          .data
		.rp_channel              (limiter_001_rsp_src_channel),                                                            //          .channel
		.rp_startofpacket        (limiter_001_rsp_src_startofpacket),                                                      //          .startofpacket
		.rp_endofpacket          (limiter_001_rsp_src_endofpacket),                                                        //          .endofpacket
		.rp_ready                (limiter_001_rsp_src_ready),                                                              //          .ready
		.av_response             (),                                                                                       // (terminated)
		.av_writeresponserequest (1'b0),                                                                                   // (terminated)
		.av_writeresponsevalid   ()                                                                                        // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_BEGIN_BURST           (90),
		.PKT_BURSTWRAP_H           (82),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BURST_SIZE_H          (85),
		.PKT_BURST_SIZE_L          (83),
		.PKT_BURST_TYPE_H          (87),
		.PKT_BURST_TYPE_L          (86),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (92),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (95),
		.PKT_THREAD_ID_H           (98),
		.PKT_THREAD_ID_L           (98),
		.PKT_CACHE_H               (105),
		.PKT_CACHE_L               (102),
		.PKT_DATA_SIDEBAND_H       (89),
		.PKT_DATA_SIDEBAND_L       (89),
		.PKT_QOS_H                 (91),
		.PKT_QOS_L                 (91),
		.PKT_ADDR_SIDEBAND_H       (88),
		.PKT_ADDR_SIDEBAND_L       (88),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_RESPONSE_STATUS_L     (106),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (5),
		.AV_BURSTCOUNT_W           (8),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) tiger_icache_icache_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                                //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.av_address              (tiger_icache_icache_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (tiger_icache_icache_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (tiger_icache_icache_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (tiger_icache_icache_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (tiger_icache_icache_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (tiger_icache_icache_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (tiger_icache_icache_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (tiger_icache_icache_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (tiger_icache_icache_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (tiger_icache_icache_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (tiger_icache_icache_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (tiger_icache_icache_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (tiger_icache_icache_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (tiger_icache_icache_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (tiger_icache_icache_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (tiger_icache_icache_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_004_src1_valid),                                                          //        rp.valid
		.rp_data                 (rsp_xbar_demux_004_src1_data),                                                           //          .data
		.rp_channel              (rsp_xbar_demux_004_src1_channel),                                                        //          .channel
		.rp_startofpacket        (rsp_xbar_demux_004_src1_startofpacket),                                                  //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_004_src1_endofpacket),                                                    //          .endofpacket
		.rp_ready                (rsp_xbar_demux_004_src1_ready),                                                          //          .ready
		.av_response             (),                                                                                       // (terminated)
		.av_writeresponserequest (1'b0),                                                                                   // (terminated)
		.av_writeresponsevalid   ()                                                                                        // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_BEGIN_BURST           (90),
		.PKT_BURSTWRAP_H           (82),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BURST_SIZE_H          (85),
		.PKT_BURST_SIZE_L          (83),
		.PKT_BURST_TYPE_H          (87),
		.PKT_BURST_TYPE_L          (86),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (92),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (95),
		.PKT_THREAD_ID_H           (98),
		.PKT_THREAD_ID_L           (98),
		.PKT_CACHE_H               (105),
		.PKT_CACHE_L               (102),
		.PKT_DATA_SIDEBAND_H       (89),
		.PKT_DATA_SIDEBAND_L       (89),
		.PKT_QOS_H                 (91),
		.PKT_QOS_L                 (91),
		.PKT_ADDR_SIDEBAND_H       (88),
		.PKT_ADDR_SIDEBAND_L       (88),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_RESPONSE_STATUS_L     (106),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (5),
		.AV_BURSTCOUNT_W           (5),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dcache_cache_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                         //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.av_address              (dcache_cache_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (dcache_cache_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (dcache_cache_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (dcache_cache_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (dcache_cache_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (dcache_cache_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (dcache_cache_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (dcache_cache_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (dcache_cache_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (dcache_cache_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (dcache_cache_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (dcache_cache_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (dcache_cache_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (dcache_cache_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (dcache_cache_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (dcache_cache_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_004_src2_valid),                                                   //        rp.valid
		.rp_data                 (rsp_xbar_demux_004_src2_data),                                                    //          .data
		.rp_channel              (rsp_xbar_demux_004_src2_channel),                                                 //          .channel
		.rp_startofpacket        (rsp_xbar_demux_004_src2_startofpacket),                                           //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_004_src2_endofpacket),                                             //          .endofpacket
		.rp_ready                (rsp_xbar_demux_004_src2_ready),                                                   //          .ready
		.av_response             (),                                                                                // (terminated)
		.av_writeresponserequest (1'b0),                                                                            // (terminated)
		.av_writeresponsevalid   ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (90),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (92),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (82),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_RESPONSE_STATUS_L     (106),
		.PKT_BURST_SIZE_H          (85),
		.PKT_BURST_SIZE_L          (83),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (108),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dcache_cache_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dcache_cache_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src0_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_src0_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_demux_src0_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_src0_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src0_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src0_channel),                                                             //                .channel
		.rf_sink_ready           (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                   //     (terminated)
		.m0_writeresponserequest (),                                                                                        //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                     //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (109),
		.FIFO_DEPTH          (5),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dcache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (90),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (92),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (82),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_RESPONSE_STATUS_L     (106),
		.PKT_BURST_SIZE_H          (85),
		.PKT_BURST_SIZE_L          (83),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (108),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                                       //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                                       //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                                        //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                                     //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (109),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (90),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (92),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (82),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_RESPONSE_STATUS_L     (106),
		.PKT_BURST_SIZE_H          (85),
		.PKT_BURST_SIZE_L          (83),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (108),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) uart_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                           //       clk_reset.reset
		.m0_address              (uart_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (uart_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (uart_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (uart_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (uart_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (uart_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (uart_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (uart_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (uart_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (uart_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (uart_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (uart_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (uart_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (uart_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (uart_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (uart_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src2_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_src2_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_src2_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_src2_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src2_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src2_channel),                                                  //                .channel
		.rf_sink_ready           (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (109),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.in_data           (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (90),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (94),
		.PKT_SRC_ID_L              (92),
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (95),
		.PKT_BURSTWRAP_H           (82),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_RESPONSE_STATUS_L     (106),
		.PKT_BURST_SIZE_H          (85),
		.PKT_BURST_SIZE_L          (83),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (108),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src1_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src1_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src1_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src1_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src1_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src1_channel),                                                                    //                .channel
		.rf_sink_ready           (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (109),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (79),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (64),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (83),
		.PKT_PROTECTION_L          (81),
		.PKT_RESPONSE_STATUS_H     (89),
		.PKT_RESPONSE_STATUS_L     (88),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (5),
		.ST_DATA_W                 (90),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                   //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                   //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                    //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                             //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                 //                .channel
		.rf_sink_ready           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (91),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                       //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (18),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                   // (terminated)
		.csr_read          (1'b0),                                                                    // (terminated)
		.csr_write         (1'b0),                                                                    // (terminated)
		.csr_readdata      (),                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                    // (terminated)
		.almost_full_data  (),                                                                        // (terminated)
		.almost_empty_data (),                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                    // (terminated)
		.out_startofpacket (),                                                                        // (terminated)
		.out_endofpacket   (),                                                                        // (terminated)
		.in_empty          (1'b0),                                                                    // (terminated)
		.out_empty         (),                                                                        // (terminated)
		.in_error          (1'b0),                                                                    // (terminated)
		.out_error         (),                                                                        // (terminated)
		.in_channel        (1'b0),                                                                    // (terminated)
		.out_channel       ()                                                                         // (terminated)
	);

	legup_system_addr_router addr_router (
		.sink_ready         (tiger_mips_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (tiger_mips_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (tiger_mips_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (tiger_mips_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (tiger_mips_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                              //       src.ready
		.src_valid          (addr_router_src_valid),                                                              //          .valid
		.src_data           (addr_router_src_data),                                                               //          .data
		.src_channel        (addr_router_src_channel),                                                            //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                         //          .endofpacket
	);

	legup_system_addr_router_001 addr_router_001 (
		.sink_ready         (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_to_fpga_bridge_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                              //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                              //          .valid
		.src_data           (addr_router_001_src_data),                                                               //          .data
		.src_channel        (addr_router_001_src_channel),                                                            //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                         //          .endofpacket
	);

	legup_system_addr_router_002 addr_router_002 (
		.sink_ready         (tiger_icache_icache_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (tiger_icache_icache_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (tiger_icache_icache_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (tiger_icache_icache_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (tiger_icache_icache_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                              //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                              //          .valid
		.src_data           (addr_router_002_src_data),                                                               //          .data
		.src_channel        (addr_router_002_src_channel),                                                            //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                         //          .endofpacket
	);

	legup_system_addr_router_002 addr_router_003 (
		.sink_ready         (dcache_cache_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (dcache_cache_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (dcache_cache_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (dcache_cache_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dcache_cache_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                       //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                       //          .valid
		.src_data           (addr_router_003_src_data),                                                        //          .data
		.src_channel        (addr_router_003_src_channel),                                                     //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                                  //          .endofpacket
	);

	legup_system_id_router id_router (
		.sink_ready         (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dcache_cache_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                           //       src.ready
		.src_valid          (id_router_src_valid),                                                           //          .valid
		.src_data           (id_router_src_data),                                                            //          .data
		.src_channel        (id_router_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                      //          .endofpacket
	);

	legup_system_id_router_001 id_router_001 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                                //       src.ready
		.src_valid          (id_router_001_src_valid),                                                                //          .valid
		.src_data           (id_router_001_src_data),                                                                 //          .data
		.src_channel        (id_router_001_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                           //          .endofpacket
	);

	legup_system_id_router id_router_002 (
		.sink_ready         (uart_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (uart_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (uart_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (uart_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (uart_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                 // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                            //       src.ready
		.src_valid          (id_router_002_src_valid),                                            //          .valid
		.src_data           (id_router_002_src_data),                                             //          .data
		.src_channel        (id_router_002_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                       //          .endofpacket
	);

	legup_system_id_router_003 id_router_003 (
		.sink_ready         (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (leap_sim_control_bridge_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_003_src_valid),                                                                  //          .valid
		.src_data           (id_router_003_src_data),                                                                   //          .data
		.src_channel        (id_router_003_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                             //          .endofpacket
	);

	legup_system_id_router_004 id_router_004 (
		.sink_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                             //       src.ready
		.src_valid          (id_router_004_src_valid),                                             //          .valid
		.src_data           (id_router_004_src_data),                                              //          .data
		.src_channel        (id_router_004_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                        //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (95),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (4),
		.PIPELINED                 (0),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (5),
		.VALID_WIDTH               (5),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clk_clk),                        //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (97),
		.PKT_DEST_ID_L             (95),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (5),
		.VALID_WIDTH               (5),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (clk_clk),                            //       clk.clk
		.reset                  (rst_controller_001_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_001_src_data),           //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (72),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.PKT_BURST_TYPE_H          (69),
		.PKT_BURST_TYPE_L          (68),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (64),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (90),
		.ST_CHANNEL_W              (5),
		.OUT_BYTE_CNT_H            (57),
		.OUT_BURSTWRAP_H           (64),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (1),
		.BURSTWRAP_CONST_VALUE     (1)
	) burst_adapter (
		.clk                   (clk_clk),                             //       cr0.clk
		.reset                 (rst_controller_001_reset_out_reset),  // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                           // reset_in0.reset
		.reset_in1  (leap_profiler_leap_processor_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                                  //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),           // reset_out.reset
		.reset_req  (),                                         // (terminated)
		.reset_in2  (1'b0),                                     // (terminated)
		.reset_in3  (1'b0),                                     // (terminated)
		.reset_in4  (1'b0),                                     // (terminated)
		.reset_in5  (1'b0),                                     // (terminated)
		.reset_in6  (1'b0),                                     // (terminated)
		.reset_in7  (1'b0),                                     // (terminated)
		.reset_in8  (1'b0),                                     // (terminated)
		.reset_in9  (1'b0),                                     // (terminated)
		.reset_in10 (1'b0),                                     // (terminated)
		.reset_in11 (1'b0),                                     // (terminated)
		.reset_in12 (1'b0),                                     // (terminated)
		.reset_in13 (1'b0),                                     // (terminated)
		.reset_in14 (1'b0),                                     // (terminated)
		.reset_in15 (1'b0)                                      // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	legup_system_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                           //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket)    //           .endofpacket
	);

	legup_system_cmd_xbar_demux cmd_xbar_demux_001 (
		.clk                (clk_clk),                               //        clk.clk
		.reset              (rst_controller_001_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_001_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_001_cmd_src_channel),           //           .channel
		.sink_data          (limiter_001_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_001_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_001_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_001_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //           .endofpacket
	);

	legup_system_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	legup_system_cmd_xbar_demux_002 cmd_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_003_src_ready),             //      sink.ready
		.sink_channel       (addr_router_003_src_channel),           //          .channel
		.sink_data          (addr_router_003_src_data),              //          .data
		.sink_startofpacket (addr_router_003_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_003_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_003_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	legup_system_cmd_xbar_mux_001 cmd_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	legup_system_cmd_xbar_mux_004 cmd_xbar_mux_004 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_004_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_004_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_004_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_004_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_004_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_004_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src2_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_003_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	legup_system_cmd_xbar_demux_002 rsp_xbar_demux (
		.clk                (clk_clk),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sink_ready         (id_router_src_ready),                //      sink.ready
		.sink_channel       (id_router_src_channel),              //          .channel
		.sink_data          (id_router_src_data),                 //          .data
		.sink_startofpacket (id_router_src_startofpacket),        //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),          //          .endofpacket
		.sink_valid         (id_router_src_valid),                //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),          //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),           //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket)     //          .endofpacket
	);

	legup_system_rsp_xbar_demux_001 rsp_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	legup_system_cmd_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	legup_system_cmd_xbar_demux_002 rsp_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	legup_system_rsp_xbar_demux_004 rsp_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_004_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_004_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_004_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_004_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_004_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_004_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_004_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_004_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_004_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_004_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_004_src2_endofpacket)    //          .endofpacket
	);

	legup_system_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	legup_system_rsp_xbar_mux rsp_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_001_src1_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_003_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_004_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (81),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (82),
		.IN_PKT_BURSTWRAP_L            (82),
		.IN_PKT_BURST_SIZE_H           (85),
		.IN_PKT_BURST_SIZE_L           (83),
		.IN_PKT_RESPONSE_STATUS_H      (107),
		.IN_PKT_RESPONSE_STATUS_L      (106),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (87),
		.IN_PKT_BURST_TYPE_L           (86),
		.IN_ST_DATA_W                  (108),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (63),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (67),
		.OUT_PKT_BURST_SIZE_L          (65),
		.OUT_PKT_RESPONSE_STATUS_H     (89),
		.OUT_PKT_RESPONSE_STATUS_L     (88),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (69),
		.OUT_PKT_BURST_TYPE_L          (68),
		.OUT_ST_DATA_W                 (90),
		.ST_CHANNEL_W                  (5),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter (
		.clk                  (clk_clk),                            //       clk.clk
		.reset                (rst_controller_001_reset_out_reset), // clk_reset.reset
		.in_valid             (cmd_xbar_mux_004_src_valid),         //      sink.valid
		.in_channel           (cmd_xbar_mux_004_src_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_mux_004_src_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_004_src_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_mux_004_src_ready),         //          .ready
		.in_data              (cmd_xbar_mux_004_src_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_src_data),             //          .data
		.out_channel          (width_adapter_src_channel),          //          .channel
		.out_valid            (width_adapter_src_valid),            //          .valid
		.out_ready            (width_adapter_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                              // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (63),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (64),
		.IN_PKT_BURSTWRAP_L            (64),
		.IN_PKT_BURST_SIZE_H           (67),
		.IN_PKT_BURST_SIZE_L           (65),
		.IN_PKT_RESPONSE_STATUS_H      (89),
		.IN_PKT_RESPONSE_STATUS_L      (88),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (69),
		.IN_PKT_BURST_TYPE_L           (68),
		.IN_ST_DATA_W                  (90),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (81),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (85),
		.OUT_PKT_BURST_SIZE_L          (83),
		.OUT_PKT_RESPONSE_STATUS_H     (107),
		.OUT_PKT_RESPONSE_STATUS_L     (106),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (87),
		.OUT_PKT_BURST_TYPE_L          (86),
		.OUT_ST_DATA_W                 (108),
		.ST_CHANNEL_W                  (5),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (1)
	) width_adapter_001 (
		.clk                  (clk_clk),                             //       clk.clk
		.reset                (rst_controller_001_reset_out_reset),  // clk_reset.reset
		.in_valid             (id_router_004_src_valid),             //      sink.valid
		.in_channel           (id_router_004_src_channel),           //          .channel
		.in_startofpacket     (id_router_004_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_004_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_004_src_ready),             //          .ready
		.in_data              (id_router_004_src_data),              //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

endmodule
