// legup_system_tb.v

// Generated using ACDS version 13.0sp1 232 at 2015.03.21.21:34:34

`timescale 1 ps / 1 ps
module legup_system_tb (
	);

	wire         legup_system_inst_clk_bfm_clk_clk;           // legup_system_inst_clk_bfm:clk -> [SDRAM_my_partner:clk, legup_system_inst:clk_clk, legup_system_inst_reset_bfm:clk]
	wire         legup_system_inst_reset_bfm_reset_reset;     // legup_system_inst_reset_bfm:reset -> legup_system_inst:reset_reset_n
	wire         legup_system_inst_uart_wire_bfm_conduit_rxd; // legup_system_inst_uart_wire_bfm:sig_rxd -> legup_system_inst:uart_wire_rxd
	wire         legup_system_inst_uart_wire_txd;             // legup_system_inst:uart_wire_txd -> legup_system_inst_uart_wire_bfm:sig_txd
	wire         legup_system_inst_sdram_wire_cs_n;           // legup_system_inst:sdram_wire_cs_n -> SDRAM_my_partner:zs_cs_n
	wire   [1:0] legup_system_inst_sdram_wire_ba;             // legup_system_inst:sdram_wire_ba -> SDRAM_my_partner:zs_ba
	wire   [1:0] legup_system_inst_sdram_wire_dqm;            // legup_system_inst:sdram_wire_dqm -> SDRAM_my_partner:zs_dqm
	wire         legup_system_inst_sdram_wire_cke;            // legup_system_inst:sdram_wire_cke -> SDRAM_my_partner:zs_cke
	wire  [11:0] legup_system_inst_sdram_wire_addr;           // legup_system_inst:sdram_wire_addr -> SDRAM_my_partner:zs_addr
	wire         legup_system_inst_sdram_wire_we_n;           // legup_system_inst:sdram_wire_we_n -> SDRAM_my_partner:zs_we_n
	wire         legup_system_inst_sdram_wire_ras_n;          // legup_system_inst:sdram_wire_ras_n -> SDRAM_my_partner:zs_ras_n
	wire         legup_system_inst_sdram_wire_cas_n;          // legup_system_inst:sdram_wire_cas_n -> SDRAM_my_partner:zs_cas_n
	wire  [15:0] sdram_my_partner_conduit_dq;                 // [] -> [SDRAM_my_partner:zs_dq, legup_system_inst:sdram_wire_dq]

	legup_system legup_system_inst (
		.clk_clk          (legup_system_inst_clk_bfm_clk_clk),           //        clk.clk
		.reset_reset_n    (legup_system_inst_reset_bfm_reset_reset),     //      reset.reset_n
		.sdram_wire_addr  (legup_system_inst_sdram_wire_addr),           // sdram_wire.addr
		.sdram_wire_ba    (legup_system_inst_sdram_wire_ba),             //           .ba
		.sdram_wire_cas_n (legup_system_inst_sdram_wire_cas_n),          //           .cas_n
		.sdram_wire_cke   (legup_system_inst_sdram_wire_cke),            //           .cke
		.sdram_wire_cs_n  (legup_system_inst_sdram_wire_cs_n),           //           .cs_n
		.sdram_wire_dq    (sdram_my_partner_conduit_dq),                 //           .dq
		.sdram_wire_dqm   (legup_system_inst_sdram_wire_dqm),            //           .dqm
		.sdram_wire_ras_n (legup_system_inst_sdram_wire_ras_n),          //           .ras_n
		.sdram_wire_we_n  (legup_system_inst_sdram_wire_we_n),           //           .we_n
		.uart_wire_rxd    (legup_system_inst_uart_wire_bfm_conduit_rxd), //  uart_wire.rxd
		.uart_wire_txd    (legup_system_inst_uart_wire_txd)              //           .txd
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) legup_system_inst_clk_bfm (
		.clk (legup_system_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) legup_system_inst_reset_bfm (
		.reset (legup_system_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (legup_system_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm legup_system_inst_uart_wire_bfm (
		.sig_rxd (legup_system_inst_uart_wire_bfm_conduit_rxd), // conduit.rxd
		.sig_txd (legup_system_inst_uart_wire_txd)              //        .txd
	);

	altera_sdram_partner_module sdram_my_partner (
		.clk      (legup_system_inst_clk_bfm_clk_clk),  //     clk.clk
		.zs_dq    (sdram_my_partner_conduit_dq),        // conduit.dq
		.zs_addr  (legup_system_inst_sdram_wire_addr),  //        .addr
		.zs_ba    (legup_system_inst_sdram_wire_ba),    //        .ba
		.zs_cas_n (legup_system_inst_sdram_wire_cas_n), //        .cas_n
		.zs_cke   (legup_system_inst_sdram_wire_cke),   //        .cke
		.zs_cs_n  (legup_system_inst_sdram_wire_cs_n),  //        .cs_n
		.zs_dqm   (legup_system_inst_sdram_wire_dqm),   //        .dqm
		.zs_ras_n (legup_system_inst_sdram_wire_ras_n), //        .ras_n
		.zs_we_n  (legup_system_inst_sdram_wire_we_n)   //        .we_n
	);

endmodule
